// **********************************************************
// * Author : 
// * Email : 
// * Create time : 
// * Last modified : 
// *
// * Filename : sram_1920x64_dp_bit_en.v
// * Description : v1.0
// * Copyright (c) : FvChip 2023. All rights reserved.
// **********************************************************
`include "define_ctrl_sram.v"

module sram_1920x64_dp_bit_en
(
    input clk_a,                          // Clock input
    input [11-1:0] addr_a,      // Group A address input
    input [64-1:0] din_a,       // Group A data input
    input ce_a,                      // Group A chip enable input (low-active)
    input wr_en_a,                      // Group A write enable input (low-active)
    input [64-1:0] bit_en_a,    // Group A bit enable input (low-active)
    output [64-1:0] dout_a, // Group A data output

    input clk_b,                          // Clock input
    input [11-1:0] addr_b,      // Group B address input
    input [64-1:0] din_b,       // Group B data input
    input ce_b,                      // Group B chip enable input (low-active)
    input wr_en_b,                      // Group B write enable input (low-active)
    input [64-1:0] bit_en_b,    // Group B bit enable input (low-active)
    output [64-1:0] dout_b  // Group B data output
);

`ifdef SRAM_MOD
    //Sram mod
    sram_mod_dp_bit_en #(
        .ADDR_WIDTH     (11), // address width parameter
        .DATA_WIDTH     (64), // data width parameter
        .ADDR_SPACE     (1920)  // address space parameter
    ) u_sram_mod_sp_bit_en
    (
        .clk_a          (clk_a      ),
        .addr_a         (addr_a     ),
        .din_a          (din_a      ),
        .ce_a           (ce_a       ),
        .wr_en_a        (wr_en_a    ),
        .bit_en_a       (bit_en_a   ),
        .dout_a         (dout_a     ),
        .clk_b          (clk_b      ),
        .addr_b         (addr_b     ),
        .din_b          (din_b      ),
        .ce_b           (ce_b       ),
        .wr_en_b        (wr_en_b    ),
        .bit_en_b       (bit_en_b   ),
        .dout_b         (dout_b     )
    );

`elsif SRAM_HL40
// `elsif SRAM_MOD
    //Sram generated by memory complier
    SRAMDP_1920x64_BE u_sramdp_1920x64_be(
        .CLKA(clk_a), 
        .QA(dout_a),
        .ADRA(addr_a), 
        .DA(din_a), 
        .WEA(~wr_en_a), 
        .WEMA(~bit_en_a), 
        .CLKB(clk_b), 
        .QB(dout_b), 
        .ADRB(addr_b), 
        .DB(64'b0), 
        .WEB(~wr_en_b), 
        .WEMB(~bit_en_b), 
        .MEA(~ce_a), 
        .MEB(~ce_b), 
        .RMEA(1'b0), 
        .RMEB(1'b0), 
        .RMA(4'b0), 
        .RMB(4'b0), 
        .LS(1'b0), 
        .TEST1A(1'b0), 
        .TEST1B(1'b0)
    );

`elsif SRAM_SMIC40
    DP_1920x32_BE u_DP_1920x32_BE_0(
        /*input           */    .CLKA     (clk_a),
        /*input           */    .CENA     (ce_a),
        /*input [a:0]     */    .AA       (addr_a),
        /*input [d:0]     */    .DA       (din_a[31:0]),
        /*input           */    .GWENA    (wr_en_a),
        /*input [d:0]     */    .WENA     (bit_en_a[31:0]),
        /*output [d:0]    */    .QA       (dout_a[31:0]),
        /*input           */    .CLKB     (clk_b),
        /*input           */    .CENB     (ce_b),
        /*input [a:0]     */    .AB       (addr_b),
        /*input [d:0]     */    .DB       (din_b[31:0]),
        /*input           */    .GWENB    (wr_en_b),
        /*input [d:0]     */    .WENB     (bit_en_b[31:0]),
        /*output [d:0]    */    .QB       (dout_b[31:0]),
        /*input [2:0]     */    .EMAA     (3'b000),
        /*input [1:0]     */    .EMAWA    (2'b00),
        /*input [2:0]     */    .EMAB     (3'b000),
        /*input [1:0]     */    .EMAWB    (2'b00),
        //test
        /*input           */    .TENA     (1'b1),
        /*input           */    .TENB     (1'b1),
        /*input           */    .RET1N    (1'b1),
        /*output          */    .CENYA    (),
        /*output [d:0]    */    .WENYA    (),
        /*output [a:0]    */    .AYA      (),
        /*output          */    .CENYB    (),
        /*output [d:0]    */    .WENYB    (),
        /*output [a:0]    */    .AYB      (),
        /*output          */    .GWENYA   (),
        /*output          */    .GWENYB   (),
        /*output [1:0]    */    .SOA      (),
        /*output [1:0]    */    .SOB      (),
        /*input           */    .TCENA    (),
        /*input [d:0]     */    .TWENA    (),
        /*input [a:0]     */    .TAA      (),
        /*input [d:0]     */    .TDA      (),
        /*input           */    .TCENB    (),
        /*input [d:0]     */    .TWENB    (),
        /*input [a:0]     */    .TAB      (),
        /*input [d:0]     */    .TDB      (),
        /*input           */    .TGWENA   (),
        /*input           */    .TGWENB   (),
        /*input [1:0]     */    .SIA      (),
        /*input           */    .SEA      (),
        /*input           */    .DFTRAMBYP(),
        /*input [1:0]     */    .SIB      (),
        /*input           */    .SEB      (),
        /*input           */    .COLLDISN ()
    );

    DP_1920x32_BE u_DP_1920x32_BE_1(
        /*input           */    .CLKA     (clk_a),
        /*input           */    .CENA     (ce_a),
        /*input [a:0]     */    .AA       (addr_a),
        /*input [d:0]     */    .DA       (din_a[63:32]),
        /*input           */    .GWENA    (wr_en_a),
        /*input [d:0]     */    .WENA     (bit_en_a[63:32]),
        /*output [d:0]    */    .QA       (dout_a[63:32]),
        /*input           */    .CLKB     (clk_b),
        /*input           */    .CENB     (ce_b),
        /*input [a:0]     */    .AB       (addr_b),
        /*input [d:0]     */    .DB       (din_b[63:32]),
        /*input           */    .GWENB    (wr_en_b),
        /*input [d:0]     */    .WENB     (bit_en_b[63:32]),
        /*output [d:0]    */    .QB       (dout_b[63:32]),
        /*input [2:0]     */    .EMAA     (3'b000),
        /*input [1:0]     */    .EMAWA    (2'b00),
        /*input [2:0]     */    .EMAB     (3'b000),
        /*input [1:0]     */    .EMAWB    (2'b00),
        //test
        /*input           */    .TENA     (1'b1),
        /*input           */    .TENB     (1'b1),
        /*input           */    .RET1N    (1'b1),
        /*output          */    .CENYA    (),
        /*output [d:0]    */    .WENYA    (),
        /*output [a:0]    */    .AYA      (),
        /*output          */    .CENYB    (),
        /*output [d:0]    */    .WENYB    (),
        /*output [a:0]    */    .AYB      (),
        /*output          */    .GWENYA   (),
        /*output          */    .GWENYB   (),
        /*output [1:0]    */    .SOA      (),
        /*output [1:0]    */    .SOB      (),
        /*input           */    .TCENA    (),
        /*input [d:0]     */    .TWENA    (),
        /*input [a:0]     */    .TAA      (),
        /*input [d:0]     */    .TDA      (),
        /*input           */    .TCENB    (),
        /*input [d:0]     */    .TWENB    (),
        /*input [a:0]     */    .TAB      (),
        /*input [d:0]     */    .TDB      (),
        /*input           */    .TGWENA   (),
        /*input           */    .TGWENB   (),
        /*input [1:0]     */    .SIA      (),
        /*input           */    .SEA      (),
        /*input           */    .DFTRAMBYP(),
        /*input [1:0]     */    .SIB      (),
        /*input           */    .SEB      (),
        /*input           */    .COLLDISN ()
    );

`endif 





endmodule