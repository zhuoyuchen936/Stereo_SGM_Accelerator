// **********************************************************
// * Author : 
// * Email : 
// * Create time : 
// * Last modified : 
// *
// * Filename : sram_270x80_dp.v
// * Description : v1.0
// * Copyright (c) : FvChip 2023. All rights reserved.
// **********************************************************
`include "define_ctrl_sram.v"

module sram_270x80_dp
(
    input clk_a,                          // Clock input
    input [9-1:0] addr_a,      // Group A address input
    input [80-1:0] din_a,       // Group A data input
    input ce_a,                      // Group A chip enable input (low-active)
    input wr_en_a,                      // Group A write enable input (low-active)
    output [80-1:0] dout_a, // Group A data output

    input clk_b,                          // Clock input
    input [9-1:0] addr_b,      // Group B address input
    input [80-1:0] din_b,       // Group B data input
    input ce_b,                      // Group B chip enable input (low-active)
    input wr_en_b,                      // Group B write enable input (low-active)
    output [80-1:0] dout_b  // Group B data output
);

`ifdef SRAM_MOD
    //Sram mod
    sram_mod_dp #(
        .ADDR_WIDTH     (9), // address width parameter
        .DATA_WIDTH     (80), // data width parameter
        .ADDR_SPACE     (270)  // address space parameter
    ) u_sram_mod_dp
    (
        .clk_a          (clk_a      ),
        .addr_a         (addr_a     ),
        .din_a          (din_a      ),
        .ce_a           (ce_a       ),
        .wr_en_a        (wr_en_a    ),
        .dout_a         (dout_a     ),
        .clk_b          (clk_b      ),
        .addr_b         (addr_b     ),
        .din_b          (din_b      ),
        .ce_b           (ce_b       ),
        .wr_en_b        (wr_en_b    ),
        .dout_b         (dout_b     )
    );

`elsif SRAM_HL40
// `elsif SRAM_MOD
    //Sram generated by memory complier
    SRAMDP_288x80 u_sramdp_288x80_be(
        .CLKA(clk_a), 
        .QA(dout_a),
        .ADRA(addr_a), 
        .DA(din_a), 
        .WEA(~wr_en_a), 
        .CLKB(clk_b), 
        .QB(dout_b), 
        .ADRB(addr_b), 
        .DB(80'b0), 
        .WEB(~wr_en_b), 
        .MEA(~ce_a), 
        .MEB(~ce_b), 
        .RMEA(1'b0), 
        .RMEB(1'b0), 
        .RMA(4'b0), 
        .RMB(4'b0), 
        .LS(1'b0), 
        .TEST1A(1'b0), 
        .TEST1B(1'b0)
    );

`elsif SRAM_SMIC40

    DP_272x80 u_DP_272x80 (
        /*input           */    .CLKA     (clk_a),
        /*input           */    .CENA     (ce_a),
        /*input [a :0]    */    .AA       (addr_a),
        /*input [d :0]    */    .DA       (din_a),
        /*input           */    .WENA     (wr_en_a),
        /*output [d :0]   */    .QA       (dout_a),
        /*input           */    .CLKB     (clk_b),
        /*input           */    .CENB     (ce_b),
        /*input [a :0]    */    .AB       (addr_b),
        /*input [d :0]    */    .DB       (din_b),
        /*input           */    .WENB     (wr_en_b),
        /*output [d :0]   */    .QB       (dout_b),
        /*input [2:0]     */    .EMAA     (3'b000),
        /*input [1:0]     */    .EMAWA    (2'b00),
        /*input [2:0]     */    .EMAB     (3'b000),
        /*input [1:0]     */    .EMAWB    (2'b00),
        //test
        /*input           */    .TENA     (1'b1),
        /*input           */    .TENB     (1'b1),
        /*input           */    .RET1N    (1'b1),
        /*output          */    .CENYA    (),
        /*output          */    .WENYA    (),
        /*output [a :0]   */    .AYA      (),
        /*output          */    .CENYB    (),
        /*output          */    .WENYB    (),
        /*output [a :0]   */    .AYB      (),
        /*output [1:0]    */    .SOA      (),
        /*output [1:0]    */    .SOB      (),
        /*input           */    .TCENA    (),
        /*input           */    .TWENA    (),
        /*input [a :0]    */    .TAA      (),
        /*input [d :0]    */    .TDA      (),
        /*input           */    .TCENB    (),
        /*input           */    .TWENB    (),
        /*input [a :0]    */    .TAB      (),
        /*input [d :0]    */    .TDB      (),
        /*input [1:0]     */    .SIA      (),
        /*input           */    .SEA      (),
        /*input           */    .DFTRAMBYP(),
        /*input [1:0]     */    .SIB      (),
        /*input           */    .SEB      (),
        /*input           */    .COLLDISN ()
    );


`endif 





endmodule