// **********************************************************
// * Author : 
// * Email : 
// * Create time : 
// * Last modified : 
// *
// * Filename : sram_2048x16_2prf.v
// * Description : v1.0
// * Copyright (c) : FvChip 2023. All rights reserved.
// **********************************************************
`include "define_ctrl_sram.v"

module sram_2048x16_2prf
(
    input clk_w,                       // Clock input
    input [11-1:0] addr_w,      // Write address input
    input [16-1:0] din_w,       // Write data input
    input ce_w,                             // Write chip enable input (low-active)
    input en_w,                             // Write enable input (low-active)
    input clk_r,                       // Clock input
    input [11-1:0] addr_r,      // Read address input
    input ce_r,                             // Read chip enable input (low-active)
    //Warning: For some memory in manufacturing processes, en_r usually not adjustable and always reading .
    input en_r,                             // Read enable input (low-active)
    output [16-1:0] dout_r  // Read data output
);

`ifdef SRAM_MOD
    //Sram mod
    sram_mod_2prf #(
        .ADDR_WIDTH     (11), // address width parameter
        .DATA_WIDTH     (16), // data width parameter
        .ADDR_SPACE     (2048)  // address space parameter
    ) u_sram_mod_2prf
    (
        .clk_w          (clk_w     ),
        .addr_w         (addr_w    ),
        .din_w          (din_w     ),
        .ce_w           (ce_w      ),
        .en_w           (en_w      ),
        .clk_r          (clk_r     ),
        .addr_r         (addr_r    ),
        .ce_r           (ce_r      ),
        .en_r           (en_r      ),
        .dout_r         (dout_r    )
    );

`elsif SRAM_HL40
// `elsif SRAM_MOD
    //Sram generated by memory complier
    SRAMDP_2048x16 u_sramdp_2048x16_be(
        .CLKA(clk_w), 
        .QA(),
        .ADRA(addr_w), 
        .DA(din_w), 
        .WEA(~en_w), 
        .CLKB(clk_r), 
        .QB(dout_r), 
        .ADRB(addr_r), 
        .DB(16'b0), 
        .WEB(~en_r), 
        .MEA(~ce_w), 
        .MEB(~ce_r), 
        .RMEA(1'b0), 
        .RMEB(1'b0), 
        .RMA(4'b0), 
        .RMB(4'b0), 
        .LS(1'b0), 
        .TADRA(11'b0), 
        .TADRB(11'b0), 
        //test port
        .DFTCLKEN(1'b0), 
        .DFTMASK(1'b0), 
        .TCLKA(1'b0), 
        .TCLKB(1'b0), 
        .BISTEA(1'b0), 
        .BISTEB(1'b0), 

        .TDA(4'b0), 
        .TWEA(1'b0), 
        .TMEA(1'b0), 
        .TCLKEA(1'b0), 
        .TEST1A(1'b0), 
        .CDA(4'b0), 
        .CAPTA(1'b0), 
        .PIPEMEA(1'b0), 
        .TPIPEMEA(1'b0), 
        .STICKYA(1'b0), 
        .SI_QA(1'b0), 
        .SI_DA(1'b0), 
        .SE_QA(1'b0), 
        .SE_INA(1'b0), 
        .SI_CNTRA(1'b0), 
        .TDB(4'b0), 
        .TWEB(1'b0), 
        .TMEB(1'b0), 
        .TCLKEB(1'b0), 
        .TEST1B(1'b0), 
        .CDB(4'b0), 
        .CAPTB(1'b0), 
        .PIPEMEB(1'b0), 
        .TPIPEMEB(1'b0), 
        .STICKYB(1'b0), 
        .SI_QB(1'b0), 
        .SI_DB(1'b0), 
        .SE_QB(1'b0), 
        .SE_INB(1'b0), 
        .SI_CNTRB(1'b0),

        .QPA(), 
        .SO_QA(), 
        .SO_DA(), 
        .SO_CNTRA(), 
        .QPB(), 
        .SO_QB(), 
        .SO_DB(), 
        .SO_CNTRB()
        
        
    );

`endif 





endmodule