module output_ABW
(
	//input
	w0,
	q1,
	D,
	A,
	B,
	temp_1,
	//output 
	output_A,
	output_B,
	output_W
);

	input [21:0] w0;
	input [2:0] q1;
	input [21:0] D;
	input [25:0] A;
	input [25:0] B;
	input [3:0] temp_1;
	output [25:0] output_A;
	output [25:0] output_B;
	output [21:0] output_W;
	
	wire [21:0] w1;
	wire [2:0] A1;
	wire [2:0] B1;
	reg [25:0] A_next;
	reg [25:0] B_next;
	
	
	assign w1= (q1 == 3'b010)?{{w0[21],w0[18:0],2'b0}-{D[20:0],1'b0}} :
	(q1 == 3'b001)?{{w0[21],w0[18:0],2'b0}-{D}}:(q1 == 3'b000)?{w0[21],w0[18:0],2'b0} :
	(q1 == 3'b111)?{{w0[21],w0[18:0],2'b0}+{D}}:{{w0[21],w0[18:0],2'b0}+{D[20:0],1'b0}};
	
	assign A1= (q1[2])?{3'b100+q1} :{3'b000};
	assign B1= (q1[2])?{3'b011+q1} :(q1==3'b000)?{3'b011+q1} :{3'b000};
	
	always@(*)
begin
    case(temp_1)
        4'd0:
        begin
		  	A_next=~q1[2]?{A[25],q1[1:0],A[22:0]}:{B[25],A1[1:0],B[22:0]};
        	B_next=~q1[2]&(|q1[1:0])?{A[25],q1[1:0]-2'b1,A[22:0]}:{B[25],B1[1:0],B[22:0]};
		 // 	A_next=~q1[2]?{A[17],q1[1:0],A[14:0]}:{B[17],A1[1:0],B[14:0]};
        	//B_next=~q1[2]&(|q1[1:0])?{A[17],q1[1:0]-2'b1,A[14:0]}:{B[17],B1[1:0],B[14:0]};
        end
        4'd1:
        begin
        	A_next=~q1[2]?{A[25:23],q1[1:0],A[20:0]}:{B[25:23],A1[1:0],B[20:0]};
        	B_next=~q1[2]&(|q1[1:0])?{A[25:23],q1[1:0]-2'b1,A[20:0]}:{B[25:23],B1[1:0],B[20:0]};
        end
		   4'd2:
        begin
        	A_next=~q1[2]?{A[25:21],q1[1:0],A[18:0]}:{B[25:21],A1[1:0],B[18:0]};
        	B_next=~q1[2]&(|q1[1:0])?{A[25:21],q1[1:0]-2'b1,A[18:0]}:{B[25:21],B1[1:0],B[18:0]};
        end
		   4'd3:
        begin
        	A_next=~q1[2]?{A[25:19],q1[1:0],A[16:0]}:{B[25:19],A1[1:0],B[16:0]};
        	B_next=~q1[2]&(|q1[1:0])?{A[25:19],q1[1:0]-2'b1,A[16:0]}:{B[25:19],B1[1:0],B[16:0]};
        end
		   4'd4:
        begin
        	A_next=~q1[2]?{A[25:17],q1[1:0],A[14:0]}:{B[25:17],A1[1:0],B[14:0]};
        	B_next=~q1[2]&(|q1[1:0])?{A[25:17],q1[1:0]-2'b1,A[14:0]}:{B[25:17],B1[1:0],B[14:0]};
        end
		  4'd5:
        begin
        	A_next=~q1[2]?{A[25:15],q1[1:0],A[12:0]}:{B[25:15],A1[1:0],B[12:0]};
        	B_next=~q1[2]&(|q1[1:0])?{A[25:15],q1[1:0]-2'b1,A[12:0]}:{B[25:15],B1[1:0],B[12:0]};
        end
		  4'd6:
        begin
        	A_next=~q1[2]?{A[25:13],q1[1:0],A[10:0]}:{B[25:13],A1[1:0],B[10:0]};
        	B_next=~q1[2]&(|q1[1:0])?{A[25:13],q1[1:0]-2'b1,A[10:0]}:{B[25:13],B1[1:0],B[10:0]};
        end
		   4'd7:
        begin
        	A_next=~q1[2]?{A[25:11],q1[1:0],A[8:0]}:{B[25:11],A1[1:0],B[8:0]};
        	B_next=~q1[2]&(|q1[1:0])?{A[25:11],q1[1:0]-2'b1,A[8:0]}:{B[25:11],B1[1:0],B[8:0]};
        end
		  4'd8:
        begin
        	A_next=~q1[2]?{A[25:9],q1[1:0],A[6:0]}:{B[25:9],A1[1:0],B[6:0]};
        	B_next=~q1[2]&(|q1[1:0])?{A[25:9],q1[1:0]-2'b1,A[6:0]}:{B[25:9],B1[1:0],B[6:0]};
        end
		  4'd9:
        begin
        	A_next=~q1[2]?{A[25:7],q1[1:0],A[4:0]}:{B[25:7],A1[1:0],B[4:0]};
        	B_next=~q1[2]&(|q1[1:0])?{A[25:7],q1[1:0]-2'b1,A[4:0]}:{B[25:7],B1[1:0],B[4:0]};
        end
		   4'd10:
        begin
        	A_next=~q1[2]?{A[25:5],q1[1:0],A[2:0]}:{B[25:5],A1[1:0],B[2:0]};
        	B_next=~q1[2]&(|q1[1:0])?{A[25:5],q1[1:0]-2'b1,A[2:0]}:{B[25:5],B1[1:0],B[2:0]};
        end
		   4'd11:
        begin
        	A_next=~q1[2]?{A[25:3],q1[1:0],A[0]}:{B[25:3],A1[1:0],B[0]};
        	B_next=~q1[2]&(|q1[1:0])?{A[25:3],q1[1:0]-2'b1,A[0]}:{B[25:3],B1[1:0],B[0]};
        end
default: 
	begin	
			A_next=26'b0;
        	B_next=26'b0;
	end
	endcase
end
	//assign A_next=~q1[2]?{A[15],q1[1:0],A[12:0]}:{B[15],A1[1:0],B[12:0]};
	//assign B_next=~q1[2]&(|q1[1:0])?{A[15],q1[1:0]-2'b1,A[12:0]}:{B[15],B1[1:0],B[12:0]};
	
	assign output_A=A_next;
	assign output_B=B_next;
	assign output_W=w1;
	
endmodule
	