// **********************************************************
// * Author : 
// * Email : 
// * Create time : 
// * Last modified : 
// *
// * Filename : sram_8192x8_2prf.v
// * Description : v1.0
// * Copyright (c) : FvChip 2023. All rights reserved.
// **********************************************************
`include "define_ctrl_sram.v"

module sram_8192x8_2prf
(
    input clk_w,                       // Clock input
    input [13-1:0] addr_w,      // Write address input
    input [8-1:0] din_w,       // Write data input
    input ce_w,                             // Write chip enable input (low-active)
    input en_w,                             // Write enable input (low-active)
    input clk_r,                       // Clock input
    input [13-1:0] addr_r,      // Read address input
    input ce_r,                             // Read chip enable input (low-active)
    //Warning: For some memory in manufacturing processes, en_r usually not adjustable and always reading .
    input en_r,                             // Read enable input (low-active)
    output [8-1:0] dout_r  // Read data output
);

`ifdef SRAM_MOD
    //Sram mod
    sram_mod_2prf #(
        .ADDR_WIDTH     (13), // address width parameter
        .DATA_WIDTH     (8), // data width parameter
        .ADDR_SPACE     (8192)  // address space parameter
    ) u_sram_mod_2prf
    (
        .clk_w          (clk_w     ),
        .addr_w         (addr_w    ),
        .din_w          (din_w     ),
        .ce_w           (ce_w      ),
        .en_w           (en_w      ),
        .clk_r          (clk_r     ),
        .addr_r         (addr_r    ),
        .ce_r           (ce_r      ),
        .en_r           (en_r      ),
        .dout_r         (dout_r    )
    );

`elsif FPGA
    //Sram generated by memory complier

   dpram_8192x8 u_dpram_8192x8 (
     .clka     (  clk_w      ),  // input wire clka
     .ena      (  1'b1          ),  // input wire ena
     .wea      ( ~en_w      ),  // input wire [0 : 0] wea
     .addra    (  addr_w     ),  // input wire [11 : 0] addra
     .dina     (  din_w     ),  // input wire [7 : 0] dina
     .clkb     (  clk_r      ),  // input wire clkb
     .enb      (  1'b1          ),  // input wire enb
     .addrb    (  addr_r     ),  // input wire [11 : 0] addrb
     .doutb    (  dout_r     )   // output wire [7 : 0] doutb
   );
`endif





endmodule
