/*
 * @Author: PingChengDong 
 * @Date: 2022-08-08 14:13:14 
 * @Last Modified by: KeLi
 * @Last Modified time: 2022-08-10 16:12:59
 */
 module DisparityMap_new(
    input  clk,
    input  rst,
    input  clken,
    input  enable,
	input  [10:0] width,
	input  [10:0] height,
    input  [8:0] range,
    input  avg_final_valid_L,
    input  avg_final_valid_R,
    input  [7:0] avgdata_L,
    input  [7:0] avgdata_R,

    input [6:0]P1,
    input [6:0]P2,
    output [15:0] disp_L,
    output [15:0] disp_R,
    output valid_final_L,
    output valid_final_R,
    /******************************************************************/
    /***************************Aggregation****************************/
    /******************************************************************/
 	output wr_en_Agg0_inst1,
    output [1151:0] BWEB_Agg0_inst1,
    output [10:0]  wr_addr_Agg0_inst1,
    output [10:0]  rd_addr_Agg0_inst1,

	input  [1151:0] Q_Aggregation0_Ram_2,
	output [1151:0] D_Aggregation0_Ram_1,

    output wr_en_Agg135_inst1,
    output [895:0] BWEB_Agg135_inst1,
    output [10:0]  wr_addr_Agg135_inst1,
    output [10:0]  rd_addr_Agg135_inst1,


	input  [895:0] Q_Aggregation135_Ram_2,
	output [895:0] D_Aggregation135_Ram_1
);
	wire   clken0 = enable | clken;

	wire [1023:0] Hamming_L;
	wire [1023:0] Hamming_R;
   	wire valid;
 	wire [7:0] disp_lrc;
	wire [6:0]disp0;
	wire valid_final_lrc;
	//census's memory
	wire  [7:0] lb0_pixel4_L;
    wire  [7:0] lb1_pixel4_L;
    wire  [7:0] lb2_pixel4_L;
    wire  [7:0] lb3_pixel4_L;

	wire  [7:0] taps0x_L;
    wire  [7:0] taps1x_L;
    wire  [7:0] taps2x_L;
    wire  [7:0] taps3x_L;
    wire  [7:0] taps4x_L;
 
    wire  [7:0] taps0x_R;
    wire  [7:0] taps1x_R;
    wire  [7:0] taps2x_R;
    wire  [7:0] taps3x_R;
    wire  [7:0] taps4x_R;

	wire [3071:0] cost_grad_R;
	wire [3071:0] cost_grad_L;
	
	census5x5_sram census5x5_sram_inst(
		.clk(clk),
    	.rst(rst),
    	.clken(clken0),
    	.width(width),
    	.avgdata_R(avgdata_R),
    	.avgdata_L(avgdata_L),
    	.avg_final_valid_R(avg_final_valid_R),
    	.avg_final_valid_L(avg_final_valid_L),
	
    	.lb0_pixel(lb0_pixel4_L),
    	.lb1_pixel(lb1_pixel4_L),
		.lb2_pixel(lb2_pixel4_L),
    	.lb3_pixel(lb3_pixel4_L),
	
    	.taps0x_L(taps0x_L),
    	.taps1x_L(taps1x_L),
    	.taps2x_L(taps2x_L),
		.taps3x_L(taps3x_L),
    	.taps4x_L(taps4x_L),

    	.taps0x_R(taps0x_R),
    	.taps1x_R(taps1x_R),
    	.taps2x_R(taps2x_R),
		.taps3x_R(taps3x_R),
    	.taps4x_R(taps4x_R)
	);

	cost_com cost_com_inst(
		.sys_clk(clk),
		.sys_rst(rst),
	//	.clken(clken0),
		.width(width),
		.clken(clken0 & avg_final_valid_L & avg_final_valid_R),

		.taps0x_L(taps0x_L),
		.taps1x_L(taps1x_L),
		.taps2x_L(taps2x_L),
		.taps3x_L(taps3x_L),
    	.taps4x_L(taps4x_L),

		.taps0x_R(taps0x_R),
		.taps1x_R(taps1x_R),
		.taps2x_R(taps2x_R),
		.taps3x_R(taps3x_R),
    	.taps4x_R(taps4x_R),
		

		.lb0_pixel6_L(lb0_pixel4_L),
		.lb1_pixel6_L(lb1_pixel4_L),
		.lb2_pixel6_L(lb2_pixel4_L),
    	.lb3_pixel6_L(lb3_pixel4_L),

		.Hamming_R(Hamming_R),
		.Hamming_L(Hamming_L),
		.cost_grad_R(cost_grad_R),
		.cost_grad_L(cost_grad_L),

		.valid(valid)
	);


	wire [1279:0]cost_fusion_L;
	wire [1279:0]cost_fusion_R;
    // cost_grad and hammingDistance fusion
	wire fusion_out_valid_L;
	wire fusion_out_valid_R;
	
	cost_fusion cost_fusion_L_inst(
		.clk(clk),
		.rst(rst),
	
		.clken(valid),
		.cost_hamming(Hamming_L),
		.cost_grad(cost_grad_L),
	
		.valid(fusion_out_valid_L),
	
		.cost_fusion(cost_fusion_L)
	);
	
	cost_fusion cost_fusion_R_inst(
		.clk(clk),
		.rst(rst),
	
		.clken(valid),
		.cost_hamming(Hamming_R),
		.cost_grad(cost_grad_R),
	
		.valid(fusion_out_valid_R),
	
		.cost_fusion(cost_fusion_R)
	);

// two census for left and right consistency detection

	wire [575:0]cost_L;
	wire [575:0]cost_R;

	wire en_L;

	wire en_R;

	jqpart1 jqpart_L(
	.rst(rst),
	.clk(clk),
	.clken(clken0),
	.valid(valid),
	
	.cost_in(cost_fusion_L),
	.cost_out(cost_L),
	
	.en(en_L)
	);
	
	jqpart1 jqpart_R(
	.rst(rst),
	.clk(clk),
	.clken(clken0),
	.valid(valid),
	
	.cost_in(cost_fusion_R),
	.cost_out(cost_R),
	
	.en(en_R)
	);
	
	reg [63:0]valid_range;
	wire [6:0] range_divide4;
	wire [8:0] range_divide4_9b;
	assign range_divide4_9b = (range>>2);
	assign range_divide4=range_divide4_9b[6:0];

	always @(*)case (range_divide4)
		7'd16: valid_range={{48{1'b0}},{16{1'b1}}};
		7'd17: valid_range={{47{1'b0}},{17{1'b1}}};
		7'd18: valid_range={{46{1'b0}},{18{1'b1}}};
		7'd19: valid_range={{45{1'b0}},{19{1'b1}}};
		7'd20: valid_range={{44{1'b0}},{20{1'b1}}};
		7'd21: valid_range={{43{1'b0}},{21{1'b1}}};
		7'd22: valid_range={{42{1'b0}},{22{1'b1}}};
		7'd23: valid_range={{41{1'b0}},{23{1'b1}}};
		7'd24: valid_range={{40{1'b0}},{24{1'b1}}};
		7'd25: valid_range={{39{1'b0}},{25{1'b1}}};
		7'd26: valid_range={{38{1'b0}},{26{1'b1}}};
		7'd27: valid_range={{37{1'b0}},{27{1'b1}}};
		7'd28: valid_range={{36{1'b0}},{28{1'b1}}};
		7'd29: valid_range={{35{1'b0}},{29{1'b1}}};
		7'd30: valid_range={{34{1'b0}},{30{1'b1}}};
		7'd31: valid_range={{33{1'b0}},{31{1'b1}}};
		7'd32: valid_range={{32{1'b0}},{32{1'b1}}};
		7'd33: valid_range={{31{1'b0}},{33{1'b1}}};
		7'd34: valid_range={{30{1'b0}},{34{1'b1}}};
		7'd35: valid_range={{29{1'b0}},{35{1'b1}}};
		7'd36: valid_range={{28{1'b0}},{36{1'b1}}};
		7'd37: valid_range={{27{1'b0}},{37{1'b1}}};
		7'd38: valid_range={{26{1'b0}},{38{1'b1}}};
		7'd39: valid_range={{25{1'b0}},{39{1'b1}}};
		7'd40: valid_range={{24{1'b0}},{40{1'b1}}};
		7'd41: valid_range={{23{1'b0}},{41{1'b1}}};
		7'd42: valid_range={{22{1'b0}},{42{1'b1}}};
		7'd43: valid_range={{21{1'b0}},{43{1'b1}}};
		7'd44: valid_range={{20{1'b0}},{44{1'b1}}};
		7'd45: valid_range={{19{1'b0}},{45{1'b1}}};
		7'd46: valid_range={{18{1'b0}},{46{1'b1}}};
		7'd47: valid_range={{17{1'b0}},{47{1'b1}}};
		7'd48: valid_range={{16{1'b0}},{48{1'b1}}};
		7'd49: valid_range={{15{1'b0}},{49{1'b1}}};
		7'd50: valid_range={{14{1'b0}},{50{1'b1}}};
		7'd51: valid_range={{13{1'b0}},{51{1'b1}}};
		7'd52: valid_range={{12{1'b0}},{52{1'b1}}};
		7'd53: valid_range={{11{1'b0}},{53{1'b1}}};
		7'd54: valid_range={{10{1'b0}},{54{1'b1}}};
		7'd55: valid_range={{9{1'b0}},{55{1'b1}}};
		7'd56: valid_range={{8{1'b0}},{56{1'b1}}};
		7'd57: valid_range={{7{1'b0}},{57{1'b1}}};
		7'd58: valid_range={{6{1'b0}},{58{1'b1}}};
		7'd59: valid_range={{5{1'b0}},{59{1'b1}}};
		7'd60: valid_range={{4{1'b0}},{60{1'b1}}};
		7'd61: valid_range={{3{1'b0}},{61{1'b1}}};
		7'd62: valid_range={{2{1'b0}},{62{1'b1}}};
		7'd63: valid_range={{1{1'b0}},{63{1'b1}}};
		7'd64: valid_range={{64{1'b1}}};
		default: valid_range={{64{1'b1}}};
	endcase


//*************************************************aggregation***************************************************************

	parameter cost_width = 9;
//connection

	wire [cost_width-1:0] cost_R_in[63:0];
	wire [cost_width-1:0] cost_L_in[63:0];
	wire [63:0] cost_valid;
	wire [(cost_width*64-1):0] cost0_valid_B;
	wire [((cost_width-2)*64-1):0] cost135_valid_B;
	assign cost_valid=valid_range;

    genvar t;
	generate for(t=0;t<64;t=t+1) begin: inloop
			// assign cost_L[t-32] = {1'd0,cost_L_temp[t-32]};
			// assign cost_R[t-32] = {1'd0,cost_R_temp[t-32]};
			assign cost_L_in[t]= cost_L[(t+1)*cost_width-1:t*cost_width] & {cost_width{valid_range[t]}};
			assign cost_R_in[t]= cost_R[(t+1)*cost_width-1:t*cost_width] & {cost_width{valid_range[t]}};
            assign cost0_valid_B[(t+1)*cost_width-1:t*cost_width] = {cost_width{~valid_range[t]}};
            assign cost135_valid_B[(t+1)*(cost_width-2)-1:t*(cost_width-2)] = {(cost_width-2){~valid_range[t]}};

		end
	endgenerate
//connection
	wire  [cost_width-1:0] min_0_R;
	
	
	reg en_first_R;
	reg en_first_R_agg2;
	wire en_agg3_R;
	
	wire [cost_width-1:0] new4_L0_R[63:0];
	wire [cost_width-3:0] new4_L135_R[63:0];
	
	
	wire  [cost_width-3:0] min_135_R;
	
	//agg3
	wire en_disp_R;
	
	wire valid_1_R;	
	wire valid_2_R;
	reg change_R;
	wire valid_3_R;
	//middle
	
	wire [cost_width-1:0] L_3_0_R[63:0];
	wire [cost_width-3:0] L_3_135_R[63:0];
	
	wire  [cost_width-1:0]L_0_R[63:0][2:0];
	wire  [cost_width-3:0]L_135_R[63:0][2:0];
	assign L_0_R[0][0]=L_3_0_R[0];
	assign L_0_R[1][0]=L_3_0_R[1];
	assign L_0_R[2][0]=L_3_0_R[2];
	assign L_0_R[3][0]=L_3_0_R[3];
	assign L_0_R[4][0]=L_3_0_R[4];
	assign L_0_R[5][0]=L_3_0_R[5];
	assign L_0_R[6][0]=L_3_0_R[6];
	assign L_0_R[7][0]=L_3_0_R[7];
	assign L_0_R[8][0]=L_3_0_R[8];
	assign L_0_R[9][0]=L_3_0_R[9];
	assign L_0_R[10][0]=L_3_0_R[10];
	assign L_0_R[11][0]=L_3_0_R[11];
	assign L_0_R[12][0]=L_3_0_R[12];
	assign L_0_R[13][0]=L_3_0_R[13];
	assign L_0_R[14][0]=L_3_0_R[14];
	assign L_0_R[15][0]=L_3_0_R[15];
	assign L_0_R[16][0]=L_3_0_R[16];
	assign L_0_R[17][0]=L_3_0_R[17];
	assign L_0_R[18][0]=L_3_0_R[18];
	assign L_0_R[19][0]=L_3_0_R[19];
	assign L_0_R[20][0]=L_3_0_R[20];
	assign L_0_R[21][0]=L_3_0_R[21];
	assign L_0_R[22][0]=L_3_0_R[22];
	assign L_0_R[23][0]=L_3_0_R[23];
	assign L_0_R[24][0]=L_3_0_R[24];
	assign L_0_R[25][0]=L_3_0_R[25];
	assign L_0_R[26][0]=L_3_0_R[26];
	assign L_0_R[27][0]=L_3_0_R[27];
	assign L_0_R[28][0]=L_3_0_R[28];
	assign L_0_R[29][0]=L_3_0_R[29];
	assign L_0_R[30][0]=L_3_0_R[30];
	assign L_0_R[31][0]=L_3_0_R[31];
	assign L_0_R[32][0]=L_3_0_R[32];
	assign L_0_R[33][0]=L_3_0_R[33];
	assign L_0_R[34][0]=L_3_0_R[34];
	assign L_0_R[35][0]=L_3_0_R[35];
	assign L_0_R[36][0]=L_3_0_R[36];
	assign L_0_R[37][0]=L_3_0_R[37];
	assign L_0_R[38][0]=L_3_0_R[38];
	assign L_0_R[39][0]=L_3_0_R[39];
	assign L_0_R[40][0]=L_3_0_R[40];
	assign L_0_R[41][0]=L_3_0_R[41];
	assign L_0_R[42][0]=L_3_0_R[42];
	assign L_0_R[43][0]=L_3_0_R[43];
	assign L_0_R[44][0]=L_3_0_R[44];
	assign L_0_R[45][0]=L_3_0_R[45];
	assign L_0_R[46][0]=L_3_0_R[46];
	assign L_0_R[47][0]=L_3_0_R[47];
	assign L_0_R[48][0]=L_3_0_R[48];
	assign L_0_R[49][0]=L_3_0_R[49];
	assign L_0_R[50][0]=L_3_0_R[50];
	assign L_0_R[51][0]=L_3_0_R[51];
	assign L_0_R[52][0]=L_3_0_R[52];
	assign L_0_R[53][0]=L_3_0_R[53];
	assign L_0_R[54][0]=L_3_0_R[54];
	assign L_0_R[55][0]=L_3_0_R[55];
	assign L_0_R[56][0]=L_3_0_R[56];
	assign L_0_R[57][0]=L_3_0_R[57];
	assign L_0_R[58][0]=L_3_0_R[58];
	assign L_0_R[59][0]=L_3_0_R[59];
	assign L_0_R[60][0]=L_3_0_R[60];
	assign L_0_R[61][0]=L_3_0_R[61];
	assign L_0_R[62][0]=L_3_0_R[62];
	assign L_0_R[63][0]=L_3_0_R[63];
	
	assign L_135_R[0][0]=L_3_135_R[0];
	assign L_135_R[1][0]=L_3_135_R[1];
	assign L_135_R[2][0]=L_3_135_R[2];
	assign L_135_R[3][0]=L_3_135_R[3];
	assign L_135_R[4][0]=L_3_135_R[4];
	assign L_135_R[5][0]=L_3_135_R[5];
	assign L_135_R[6][0]=L_3_135_R[6];
	assign L_135_R[7][0]=L_3_135_R[7];
	assign L_135_R[8][0]=L_3_135_R[8];
	assign L_135_R[9][0]=L_3_135_R[9];
	assign L_135_R[10][0]=L_3_135_R[10];
	assign L_135_R[11][0]=L_3_135_R[11];
	assign L_135_R[12][0]=L_3_135_R[12];
	assign L_135_R[13][0]=L_3_135_R[13];
	assign L_135_R[14][0]=L_3_135_R[14];
	assign L_135_R[15][0]=L_3_135_R[15];
	assign L_135_R[16][0]=L_3_135_R[16];
	assign L_135_R[17][0]=L_3_135_R[17];
	assign L_135_R[18][0]=L_3_135_R[18];
	assign L_135_R[19][0]=L_3_135_R[19];
	assign L_135_R[20][0]=L_3_135_R[20];
	assign L_135_R[21][0]=L_3_135_R[21];
	assign L_135_R[22][0]=L_3_135_R[22];
	assign L_135_R[23][0]=L_3_135_R[23];
	assign L_135_R[24][0]=L_3_135_R[24];
	assign L_135_R[25][0]=L_3_135_R[25];
	assign L_135_R[26][0]=L_3_135_R[26];
	assign L_135_R[27][0]=L_3_135_R[27];
	assign L_135_R[28][0]=L_3_135_R[28];
	assign L_135_R[29][0]=L_3_135_R[29];
	assign L_135_R[30][0]=L_3_135_R[30];
	assign L_135_R[31][0]=L_3_135_R[31];
	assign L_135_R[32][0]=L_3_135_R[32];
	assign L_135_R[33][0]=L_3_135_R[33];
	assign L_135_R[34][0]=L_3_135_R[34];
	assign L_135_R[35][0]=L_3_135_R[35];
	assign L_135_R[36][0]=L_3_135_R[36];
	assign L_135_R[37][0]=L_3_135_R[37];
	assign L_135_R[38][0]=L_3_135_R[38];
	assign L_135_R[39][0]=L_3_135_R[39];
	assign L_135_R[40][0]=L_3_135_R[40];
	assign L_135_R[41][0]=L_3_135_R[41];
	assign L_135_R[42][0]=L_3_135_R[42];
	assign L_135_R[43][0]=L_3_135_R[43];
	assign L_135_R[44][0]=L_3_135_R[44];
	assign L_135_R[45][0]=L_3_135_R[45];
	assign L_135_R[46][0]=L_3_135_R[46];
	assign L_135_R[47][0]=L_3_135_R[47];
	assign L_135_R[48][0]=L_3_135_R[48];
	assign L_135_R[49][0]=L_3_135_R[49];
	assign L_135_R[50][0]=L_3_135_R[50];
	assign L_135_R[51][0]=L_3_135_R[51];
	assign L_135_R[52][0]=L_3_135_R[52];
	assign L_135_R[53][0]=L_3_135_R[53];
	assign L_135_R[54][0]=L_3_135_R[54];
	assign L_135_R[55][0]=L_3_135_R[55];
	assign L_135_R[56][0]=L_3_135_R[56];
	assign L_135_R[57][0]=L_3_135_R[57];
	assign L_135_R[58][0]=L_3_135_R[58];
	assign L_135_R[59][0]=L_3_135_R[59];
	assign L_135_R[60][0]=L_3_135_R[60];
	assign L_135_R[61][0]=L_3_135_R[61];
	assign L_135_R[62][0]=L_3_135_R[62];
	assign L_135_R[63][0]=L_3_135_R[63];
	reg en_agg4_R;
	reg rst0_R;	
		
	
	wire [cost_width-1:0] L0_R[63:0];
	wire [cost_width-3:0] L135_R[63:0];
	agg_first#(cost_width) agg_first_right(
		.clk(clk),
		.rst(rst),
		.clken(clken0),
		.valid(en_R),
		.valid_1(valid_1_R),
		
		.cost0_0(cost_R_in[0]),
		.cost0_1(cost_R_in[1]),
		.cost0_2(cost_R_in[2]),
		.cost0_3(cost_R_in[3]),
		.cost0_4(cost_R_in[4]),
		.cost0_5(cost_R_in[5]),
		.cost0_6(cost_R_in[6]),
		.cost0_7(cost_R_in[7]),
		.cost0_8(cost_R_in[8]),
		.cost0_9(cost_R_in[9]),
		.cost0_10(cost_R_in[10]),
		.cost0_11(cost_R_in[11]),
		.cost0_12(cost_R_in[12]),
		.cost0_13(cost_R_in[13]),
		.cost0_14(cost_R_in[14]),
		.cost0_15(cost_R_in[15]),
		.cost0_16(cost_R_in[16]),
		.cost0_17(cost_R_in[17]),
		.cost0_18(cost_R_in[18]),
		.cost0_19(cost_R_in[19]),
		.cost0_20(cost_R_in[20]),
		.cost0_21(cost_R_in[21]),
		.cost0_22(cost_R_in[22]),
		.cost0_23(cost_R_in[23]),
		.cost0_24(cost_R_in[24]),
		.cost0_25(cost_R_in[25]),
		.cost0_26(cost_R_in[26]),
		.cost0_27(cost_R_in[27]),
		.cost0_28(cost_R_in[28]),
		.cost0_29(cost_R_in[29]),
		.cost0_30(cost_R_in[30]),
		.cost0_31(cost_R_in[31]),
	
		.cost0_32(cost_R_in[32]),
		.cost0_33(cost_R_in[33]),
		.cost0_34(cost_R_in[34]),
		.cost0_35(cost_R_in[35]),
		.cost0_36(cost_R_in[36]),
		.cost0_37(cost_R_in[37]),
		.cost0_38(cost_R_in[38]),
		.cost0_39(cost_R_in[39]),
		.cost0_40(cost_R_in[40]),
		.cost0_41(cost_R_in[41]),
		.cost0_42(cost_R_in[42]),
		.cost0_43(cost_R_in[43]),
		.cost0_44(cost_R_in[44]),
		.cost0_45(cost_R_in[45]),
		.cost0_46(cost_R_in[46]),
		.cost0_47(cost_R_in[47]),
		.cost0_48(cost_R_in[48]),
		.cost0_49(cost_R_in[49]),
		.cost0_50(cost_R_in[50]),
		.cost0_51(cost_R_in[51]),
		.cost0_52(cost_R_in[52]),
		.cost0_53(cost_R_in[53]),
		.cost0_54(cost_R_in[54]),
		.cost0_55(cost_R_in[55]),
		.cost0_56(cost_R_in[56]),
		.cost0_57(cost_R_in[57]),
		.cost0_58(cost_R_in[58]),
		.cost0_59(cost_R_in[59]),
		.cost0_60(cost_R_in[60]),
		.cost0_61(cost_R_in[61]),
		.cost0_62(cost_R_in[62]),
		.cost0_63(cost_R_in[63]),
		
		.cost135_0(cost_R_in[0][cost_width-1:2]),
		.cost135_1(cost_R_in[1][cost_width-1:2]),
		.cost135_2(cost_R_in[2][cost_width-1:2]),
		.cost135_3(cost_R_in[3][cost_width-1:2]),
		.cost135_4(cost_R_in[4][cost_width-1:2]),
		.cost135_5(cost_R_in[5][cost_width-1:2]),
		.cost135_6(cost_R_in[6][cost_width-1:2]),
		.cost135_7(cost_R_in[7][cost_width-1:2]),
		.cost135_8(cost_R_in[8][cost_width-1:2]),
		.cost135_9(cost_R_in[9][cost_width-1:2]),
		.cost135_10(cost_R_in[10][cost_width-1:2]),
		.cost135_11(cost_R_in[11][cost_width-1:2]),
		.cost135_12(cost_R_in[12][cost_width-1:2]),
		.cost135_13(cost_R_in[13][cost_width-1:2]),
		.cost135_14(cost_R_in[14][cost_width-1:2]),
		.cost135_15(cost_R_in[15][cost_width-1:2]),
		.cost135_16(cost_R_in[16][cost_width-1:2]),
		.cost135_17(cost_R_in[17][cost_width-1:2]),
		.cost135_18(cost_R_in[18][cost_width-1:2]),
		.cost135_19(cost_R_in[19][cost_width-1:2]),
		.cost135_20(cost_R_in[20][cost_width-1:2]),
		.cost135_21(cost_R_in[21][cost_width-1:2]),
		.cost135_22(cost_R_in[22][cost_width-1:2]),
		.cost135_23(cost_R_in[23][cost_width-1:2]),
		.cost135_24(cost_R_in[24][cost_width-1:2]),
		.cost135_25(cost_R_in[25][cost_width-1:2]),
		.cost135_26(cost_R_in[26][cost_width-1:2]),
		.cost135_27(cost_R_in[27][cost_width-1:2]),
		.cost135_28(cost_R_in[28][cost_width-1:2]),
		.cost135_29(cost_R_in[29][cost_width-1:2]),
		.cost135_30(cost_R_in[30][cost_width-1:2]),
		.cost135_31(cost_R_in[31][cost_width-1:2]),
	
		.cost135_32(cost_R_in[32][cost_width-1:2]),
		.cost135_33(cost_R_in[33][cost_width-1:2]),
		.cost135_34(cost_R_in[34][cost_width-1:2]),
		.cost135_35(cost_R_in[35][cost_width-1:2]),
		.cost135_36(cost_R_in[36][cost_width-1:2]),
		.cost135_37(cost_R_in[37][cost_width-1:2]),
		.cost135_38(cost_R_in[38][cost_width-1:2]),
		.cost135_39(cost_R_in[39][cost_width-1:2]),
		.cost135_40(cost_R_in[40][cost_width-1:2]),
		.cost135_41(cost_R_in[41][cost_width-1:2]),
		.cost135_42(cost_R_in[42][cost_width-1:2]),
		.cost135_43(cost_R_in[43][cost_width-1:2]),
		.cost135_44(cost_R_in[44][cost_width-1:2]),
		.cost135_45(cost_R_in[45][cost_width-1:2]),
		.cost135_46(cost_R_in[46][cost_width-1:2]),
		.cost135_47(cost_R_in[47][cost_width-1:2]),
		.cost135_48(cost_R_in[48][cost_width-1:2]),
		.cost135_49(cost_R_in[49][cost_width-1:2]),
		.cost135_50(cost_R_in[50][cost_width-1:2]),
		.cost135_51(cost_R_in[51][cost_width-1:2]),
		.cost135_52(cost_R_in[52][cost_width-1:2]),
		.cost135_53(cost_R_in[53][cost_width-1:2]),
		.cost135_54(cost_R_in[54][cost_width-1:2]),
		.cost135_55(cost_R_in[55][cost_width-1:2]),
		.cost135_56(cost_R_in[56][cost_width-1:2]),
		.cost135_57(cost_R_in[57][cost_width-1:2]),
		.cost135_58(cost_R_in[58][cost_width-1:2]),
		.cost135_59(cost_R_in[59][cost_width-1:2]),
		.cost135_60(cost_R_in[60][cost_width-1:2]),
		.cost135_61(cost_R_in[61][cost_width-1:2]),
		.cost135_62(cost_R_in[62][cost_width-1:2]),
		.cost135_63(cost_R_in[63][cost_width-1:2]),
		
		.L0_0(L0_R[0]),
		.L0_1(L0_R[1]),
		.L0_2(L0_R[2]),
		.L0_3(L0_R[3]),
		.L0_4(L0_R[4]),
		.L0_5(L0_R[5]),
		.L0_6(L0_R[6]),
		.L0_7(L0_R[7]),
		.L0_8(L0_R[8]),
		.L0_9(L0_R[9]),
		.L0_10(L0_R[10]),
		.L0_11(L0_R[11]),
		.L0_12(L0_R[12]),
		.L0_13(L0_R[13]),
		.L0_14(L0_R[14]),
		.L0_15(L0_R[15]),
		.L0_16(L0_R[16]),
		.L0_17(L0_R[17]),
		.L0_18(L0_R[18]),
		.L0_19(L0_R[19]),
		.L0_20(L0_R[20]),
		.L0_21(L0_R[21]),
		.L0_22(L0_R[22]),
		.L0_23(L0_R[23]),
		.L0_24(L0_R[24]),
		.L0_25(L0_R[25]),
		.L0_26(L0_R[26]),
		.L0_27(L0_R[27]),
		.L0_28(L0_R[28]),
		.L0_29(L0_R[29]),
		.L0_30(L0_R[30]),
		.L0_31(L0_R[31]),
	
		.L0_32(L0_R[32]),
		.L0_33(L0_R[33]),
		.L0_34(L0_R[34]),
		.L0_35(L0_R[35]),
		.L0_36(L0_R[36]),
		.L0_37(L0_R[37]),
		.L0_38(L0_R[38]),
		.L0_39(L0_R[39]),
		.L0_40(L0_R[40]),
		.L0_41(L0_R[41]),
		.L0_42(L0_R[42]),
		.L0_43(L0_R[43]),
		.L0_44(L0_R[44]),
		.L0_45(L0_R[45]),
		.L0_46(L0_R[46]),
		.L0_47(L0_R[47]),
		.L0_48(L0_R[48]),
		.L0_49(L0_R[49]),
		.L0_50(L0_R[50]),
		.L0_51(L0_R[51]),
		.L0_52(L0_R[52]),
		.L0_53(L0_R[53]),
		.L0_54(L0_R[54]),
		.L0_55(L0_R[55]),
		.L0_56(L0_R[56]),
		.L0_57(L0_R[57]),
		.L0_58(L0_R[58]),
		.L0_59(L0_R[59]),
		.L0_60(L0_R[60]),
		.L0_61(L0_R[61]),
		.L0_62(L0_R[62]),
		.L0_63(L0_R[63]),
		
		.L135_0(L135_R[0]),
		.L135_1(L135_R[1]),
		.L135_2(L135_R[2]),
		.L135_3(L135_R[3]),
		.L135_4(L135_R[4]),
		.L135_5(L135_R[5]),
		.L135_6(L135_R[6]),
		.L135_7(L135_R[7]),
		.L135_8(L135_R[8]),
		.L135_9(L135_R[9]),
		.L135_10(L135_R[10]),
		.L135_11(L135_R[11]),
		.L135_12(L135_R[12]),
		.L135_13(L135_R[13]),
		.L135_14(L135_R[14]),
		.L135_15(L135_R[15]),
		.L135_16(L135_R[16]),
		.L135_17(L135_R[17]),
		.L135_18(L135_R[18]),
		.L135_19(L135_R[19]),
		.L135_20(L135_R[20]),
		.L135_21(L135_R[21]),
		.L135_22(L135_R[22]),
		.L135_23(L135_R[23]),
		.L135_24(L135_R[24]),
		.L135_25(L135_R[25]),
		.L135_26(L135_R[26]),
		.L135_27(L135_R[27]),
		.L135_28(L135_R[28]),
		.L135_29(L135_R[29]),
		.L135_30(L135_R[30]),
		.L135_31(L135_R[31]),
	
		.L135_32(L135_R[32]),
		.L135_33(L135_R[33]),
		.L135_34(L135_R[34]),
		.L135_35(L135_R[35]),
		.L135_36(L135_R[36]),
		.L135_37(L135_R[37]),
		.L135_38(L135_R[38]),
		.L135_39(L135_R[39]),
		.L135_40(L135_R[40]),
		.L135_41(L135_R[41]),
		.L135_42(L135_R[42]),
		.L135_43(L135_R[43]),
		.L135_44(L135_R[44]),
		.L135_45(L135_R[45]),
		.L135_46(L135_R[46]),
		.L135_47(L135_R[47]),
		.L135_48(L135_R[48]),
		.L135_49(L135_R[49]),
		.L135_50(L135_R[50]),
		.L135_51(L135_R[51]),
		.L135_52(L135_R[52]),
		.L135_53(L135_R[53]),
		.L135_54(L135_R[54]),
		.L135_55(L135_R[55]),
		.L135_56(L135_R[56]),
		.L135_57(L135_R[57]),
		.L135_58(L135_R[58]),
		.L135_59(L135_R[59]),
		.L135_60(L135_R[60]),
		.L135_61(L135_R[61]),
		.L135_62(L135_R[62]),
		.L135_63(L135_R[63])
		);
	
	wire [cost_width-1:0] L_2_0_R   [63:0];
	wire [cost_width-3:0] L_2_135_R [63:0];
	
	agg_second#(cost_width) agg_second_right(
		.clk(clk),
		.rst(rst),
		.clken(clken0),
		.valid_1(valid_1_R),
		.valid_2(valid_2_R),
		.cost0_0(L0_R[0]),
		.cost0_1(L0_R[1]),
		.cost0_2(L0_R[2]),
		.cost0_3(L0_R[3]),
		.cost0_4(L0_R[4]),
		.cost0_5(L0_R[5]),
		.cost0_6(L0_R[6]),
		.cost0_7(L0_R[7]),
		.cost0_8(L0_R[8]),
		.cost0_9(L0_R[9]),
		.cost0_10(L0_R[10]),
		.cost0_11(L0_R[11]),
		.cost0_12(L0_R[12]),
		.cost0_13(L0_R[13]),
		.cost0_14(L0_R[14]),
		.cost0_15(L0_R[15]),
		.cost0_16(L0_R[16]),
		.cost0_17(L0_R[17]),
		.cost0_18(L0_R[18]),
		.cost0_19(L0_R[19]),
		.cost0_20(L0_R[20]),
		.cost0_21(L0_R[21]),
		.cost0_22(L0_R[22]),
		.cost0_23(L0_R[23]),
		.cost0_24(L0_R[24]),
		.cost0_25(L0_R[25]),
		.cost0_26(L0_R[26]),
		.cost0_27(L0_R[27]),
		.cost0_28(L0_R[28]),
		.cost0_29(L0_R[29]),
		.cost0_30(L0_R[30]),
		.cost0_31(L0_R[31]),
		.cost0_32(L0_R[32]),
		.cost0_33(L0_R[33]),
		.cost0_34(L0_R[34]),
		.cost0_35(L0_R[35]),
		.cost0_36(L0_R[36]),
		.cost0_37(L0_R[37]),
		.cost0_38(L0_R[38]),
		.cost0_39(L0_R[39]),
		.cost0_40(L0_R[40]),
		.cost0_41(L0_R[41]),
		.cost0_42(L0_R[42]),
		.cost0_43(L0_R[43]),
		.cost0_44(L0_R[44]),
		.cost0_45(L0_R[45]),
		.cost0_46(L0_R[46]),
		.cost0_47(L0_R[47]),
		.cost0_48(L0_R[48]),
		.cost0_49(L0_R[49]),
		.cost0_50(L0_R[50]),
		.cost0_51(L0_R[51]),
		.cost0_52(L0_R[52]),
		.cost0_53(L0_R[53]),
		.cost0_54(L0_R[54]),
		.cost0_55(L0_R[55]),
		.cost0_56(L0_R[56]),
		.cost0_57(L0_R[57]),
		.cost0_58(L0_R[58]),
		.cost0_59(L0_R[59]),
		.cost0_60(L0_R[60]),
		.cost0_61(L0_R[61]),
		.cost0_62(L0_R[62]),
		.cost0_63(L0_R[63]),
	
		.cost135_0(L135_R[0]),
		.cost135_1(L135_R[1]),
		.cost135_2(L135_R[2]),
		.cost135_3(L135_R[3]),
		.cost135_4(L135_R[4]),
		.cost135_5(L135_R[5]),
		.cost135_6(L135_R[6]),
		.cost135_7(L135_R[7]),
		.cost135_8(L135_R[8]),
		.cost135_9(L135_R[9]),
		.cost135_10(L135_R[10]),
		.cost135_11(L135_R[11]),
		.cost135_12(L135_R[12]),
		.cost135_13(L135_R[13]),
		.cost135_14(L135_R[14]),
		.cost135_15(L135_R[15]),
		.cost135_16(L135_R[16]),
		.cost135_17(L135_R[17]),
		.cost135_18(L135_R[18]),
		.cost135_19(L135_R[19]),
		.cost135_20(L135_R[20]),
		.cost135_21(L135_R[21]),
		.cost135_22(L135_R[22]),
		.cost135_23(L135_R[23]),
		.cost135_24(L135_R[24]),
		.cost135_25(L135_R[25]),
		.cost135_26(L135_R[26]),
		.cost135_27(L135_R[27]),
		.cost135_28(L135_R[28]),
		.cost135_29(L135_R[29]),
		.cost135_30(L135_R[30]),
		.cost135_31(L135_R[31]),
		.cost135_32(L135_R[32]),
		.cost135_33(L135_R[33]),
		.cost135_34(L135_R[34]),
		.cost135_35(L135_R[35]),
		.cost135_36(L135_R[36]),
		.cost135_37(L135_R[37]),
		.cost135_38(L135_R[38]),
		.cost135_39(L135_R[39]),
		.cost135_40(L135_R[40]),
		.cost135_41(L135_R[41]),
		.cost135_42(L135_R[42]),
		.cost135_43(L135_R[43]),
		.cost135_44(L135_R[44]),
		.cost135_45(L135_R[45]),
		.cost135_46(L135_R[46]),
		.cost135_47(L135_R[47]),
		.cost135_48(L135_R[48]),
		.cost135_49(L135_R[49]),
		.cost135_50(L135_R[50]),
		.cost135_51(L135_R[51]),
		.cost135_52(L135_R[52]),
		.cost135_53(L135_R[53]),
		.cost135_54(L135_R[54]),
		.cost135_55(L135_R[55]),
		.cost135_56(L135_R[56]),
		.cost135_57(L135_R[57]),
		.cost135_58(L135_R[58]),
		.cost135_59(L135_R[59]),
		.cost135_60(L135_R[60]),
		.cost135_61(L135_R[61]),
		.cost135_62(L135_R[62]),
		.cost135_63(L135_R[63]),
		
		
		.L0_0(L_2_0_R[0]),
		.L0_1(L_2_0_R[1]),
		.L0_2(L_2_0_R[2]),
		.L0_3(L_2_0_R[3]),
		.L0_4(L_2_0_R[4]),
		.L0_5(L_2_0_R[5]),
		.L0_6(L_2_0_R[6]),
		.L0_7(L_2_0_R[7]),
		.L0_8(L_2_0_R[8]),
		.L0_9(L_2_0_R[9]),
		.L0_10(L_2_0_R[10]),
		.L0_11(L_2_0_R[11]),
		.L0_12(L_2_0_R[12]),
		.L0_13(L_2_0_R[13]),
		.L0_14(L_2_0_R[14]),
		.L0_15(L_2_0_R[15]),
		.L0_16(L_2_0_R[16]),
		.L0_17(L_2_0_R[17]),
		.L0_18(L_2_0_R[18]),
		.L0_19(L_2_0_R[19]),
		.L0_20(L_2_0_R[20]),
		.L0_21(L_2_0_R[21]),
		.L0_22(L_2_0_R[22]),
		.L0_23(L_2_0_R[23]),
		.L0_24(L_2_0_R[24]),
		.L0_25(L_2_0_R[25]),
		.L0_26(L_2_0_R[26]),
		.L0_27(L_2_0_R[27]),
		.L0_28(L_2_0_R[28]),
		.L0_29(L_2_0_R[29]),
		.L0_30(L_2_0_R[30]),
		.L0_31(L_2_0_R[31]),
		.L0_32(L_2_0_R[32]),
		.L0_33(L_2_0_R[33]),
		.L0_34(L_2_0_R[34]),
		.L0_35(L_2_0_R[35]),
		.L0_36(L_2_0_R[36]),
		.L0_37(L_2_0_R[37]),
		.L0_38(L_2_0_R[38]),
		.L0_39(L_2_0_R[39]),
		.L0_40(L_2_0_R[40]),
		.L0_41(L_2_0_R[41]),
		.L0_42(L_2_0_R[42]),
		.L0_43(L_2_0_R[43]),
		.L0_44(L_2_0_R[44]),
		.L0_45(L_2_0_R[45]),
		.L0_46(L_2_0_R[46]),
		.L0_47(L_2_0_R[47]),
		.L0_48(L_2_0_R[48]),
		.L0_49(L_2_0_R[49]),
		.L0_50(L_2_0_R[50]),
		.L0_51(L_2_0_R[51]),
		.L0_52(L_2_0_R[52]),
		.L0_53(L_2_0_R[53]),
		.L0_54(L_2_0_R[54]),
		.L0_55(L_2_0_R[55]),
		.L0_56(L_2_0_R[56]),
		.L0_57(L_2_0_R[57]),
		.L0_58(L_2_0_R[58]),
		.L0_59(L_2_0_R[59]),
		.L0_60(L_2_0_R[60]),
		.L0_61(L_2_0_R[61]),
		.L0_62(L_2_0_R[62]),
		.L0_63(L_2_0_R[63]),	
		
		.L135_0(L_2_135_R[0]),
		.L135_1(L_2_135_R[1]),
		.L135_2(L_2_135_R[2]),
		.L135_3(L_2_135_R[3]),
		.L135_4(L_2_135_R[4]),
		.L135_5(L_2_135_R[5]),
		.L135_6(L_2_135_R[6]),
		.L135_7(L_2_135_R[7]),
		.L135_8(L_2_135_R[8]),
		.L135_9(L_2_135_R[9]),
		.L135_10(L_2_135_R[10]),
		.L135_11(L_2_135_R[11]),
		.L135_12(L_2_135_R[12]),
		.L135_13(L_2_135_R[13]),
		.L135_14(L_2_135_R[14]),
		.L135_15(L_2_135_R[15]),
		.L135_16(L_2_135_R[16]),
		.L135_17(L_2_135_R[17]),
		.L135_18(L_2_135_R[18]),
		.L135_19(L_2_135_R[19]),
		.L135_20(L_2_135_R[20]),
		.L135_21(L_2_135_R[21]),
		.L135_22(L_2_135_R[22]),
		.L135_23(L_2_135_R[23]),
		.L135_24(L_2_135_R[24]),
		.L135_25(L_2_135_R[25]),
		.L135_26(L_2_135_R[26]),
		.L135_27(L_2_135_R[27]),
		.L135_28(L_2_135_R[28]),
		.L135_29(L_2_135_R[29]),
		.L135_30(L_2_135_R[30]),
		.L135_31(L_2_135_R[31]),
		.L135_32(L_2_135_R[32]),
		.L135_33(L_2_135_R[33]),
		.L135_34(L_2_135_R[34]),
		.L135_35(L_2_135_R[35]),
		.L135_36(L_2_135_R[36]),
		.L135_37(L_2_135_R[37]),
		.L135_38(L_2_135_R[38]),
		.L135_39(L_2_135_R[39]),
		.L135_40(L_2_135_R[40]),
		.L135_41(L_2_135_R[41]),
		.L135_42(L_2_135_R[42]),
		.L135_43(L_2_135_R[43]),
		.L135_44(L_2_135_R[44]),
		.L135_45(L_2_135_R[45]),
		.L135_46(L_2_135_R[46]),
		.L135_47(L_2_135_R[47]),
		.L135_48(L_2_135_R[48]),
		.L135_49(L_2_135_R[49]),
		.L135_50(L_2_135_R[50]),
		.L135_51(L_2_135_R[51]),
		.L135_52(L_2_135_R[52]),
		.L135_53(L_2_135_R[53]),
		.L135_54(L_2_135_R[54]),
		.L135_55(L_2_135_R[55]),
		.L135_56(L_2_135_R[56]),
		.L135_57(L_2_135_R[57]),
		.L135_58(L_2_135_R[58]),
		.L135_59(L_2_135_R[59]),
		.L135_60(L_2_135_R[60]),
		.L135_61(L_2_135_R[61]),
		.L135_62(L_2_135_R[62]),
		.L135_63(L_2_135_R[63])
	
		);
	
	wire [cost_width-1:0] new3_L0_R[63:0];
	wire [cost_width-3:0] new3_L135_R[63:0];
	
	third_agg#(cost_width) third_agg_Right(
		.clk(clk),
		.rst(rst),
		.clken(clken0),
		.change(change_R),
		.valid_2(valid_2_R),
		.valid_3(valid_3_R),
		.cost0_0(L_2_0_R[0]),
		.cost0_1(L_2_0_R[1]),
		.cost0_2(L_2_0_R[2]),
		.cost0_3(L_2_0_R[3]),
		.cost0_4(L_2_0_R[4]),
		.cost0_5(L_2_0_R[5]),
		.cost0_6(L_2_0_R[6]),
		.cost0_7(L_2_0_R[7]),
		.cost0_8(L_2_0_R[8]),
		.cost0_9(L_2_0_R[9]),
		.cost0_10(L_2_0_R[10]),
		.cost0_11(L_2_0_R[11]),
		.cost0_12(L_2_0_R[12]),
		.cost0_13(L_2_0_R[13]),
		.cost0_14(L_2_0_R[14]),
		.cost0_15(L_2_0_R[15]),
		.cost0_16(L_2_0_R[16]),
		.cost0_17(L_2_0_R[17]),
		.cost0_18(L_2_0_R[18]),
		.cost0_19(L_2_0_R[19]),
		.cost0_20(L_2_0_R[20]),
		.cost0_21(L_2_0_R[21]),
		.cost0_22(L_2_0_R[22]),
		.cost0_23(L_2_0_R[23]),
		.cost0_24(L_2_0_R[24]),
		.cost0_25(L_2_0_R[25]),
		.cost0_26(L_2_0_R[26]),
		.cost0_27(L_2_0_R[27]),
		.cost0_28(L_2_0_R[28]),
		.cost0_29(L_2_0_R[29]),
		.cost0_30(L_2_0_R[30]),
		.cost0_31(L_2_0_R[31]),
		.cost0_32(L_2_0_R[32]),
		.cost0_33(L_2_0_R[33]),
		.cost0_34(L_2_0_R[34]),
		.cost0_35(L_2_0_R[35]),
		.cost0_36(L_2_0_R[36]),
		.cost0_37(L_2_0_R[37]),
		.cost0_38(L_2_0_R[38]),
		.cost0_39(L_2_0_R[39]),
		.cost0_40(L_2_0_R[40]),
		.cost0_41(L_2_0_R[41]),
		.cost0_42(L_2_0_R[42]),
		.cost0_43(L_2_0_R[43]),
		.cost0_44(L_2_0_R[44]),
		.cost0_45(L_2_0_R[45]),
		.cost0_46(L_2_0_R[46]),
		.cost0_47(L_2_0_R[47]),
		.cost0_48(L_2_0_R[48]),
		.cost0_49(L_2_0_R[49]),
		.cost0_50(L_2_0_R[50]),
		.cost0_51(L_2_0_R[51]),
		.cost0_52(L_2_0_R[52]),
		.cost0_53(L_2_0_R[53]),
		.cost0_54(L_2_0_R[54]),
		.cost0_55(L_2_0_R[55]),
		.cost0_56(L_2_0_R[56]),
		.cost0_57(L_2_0_R[57]),
		.cost0_58(L_2_0_R[58]),
		.cost0_59(L_2_0_R[59]),
		.cost0_60(L_2_0_R[60]),
		.cost0_61(L_2_0_R[61]),
		.cost0_62(L_2_0_R[62]),
		.cost0_63(L_2_0_R[63]),
	
		.cost135_0(L_2_135_R[0]),
		.cost135_1(L_2_135_R[1]),
		.cost135_2(L_2_135_R[2]),
		.cost135_3(L_2_135_R[3]),
		.cost135_4(L_2_135_R[4]),
		.cost135_5(L_2_135_R[5]),
		.cost135_6(L_2_135_R[6]),
		.cost135_7(L_2_135_R[7]),
		.cost135_8(L_2_135_R[8]),
		.cost135_9(L_2_135_R[9]),
		.cost135_10(L_2_135_R[10]),
		.cost135_11(L_2_135_R[11]),
		.cost135_12(L_2_135_R[12]),
		.cost135_13(L_2_135_R[13]),
		.cost135_14(L_2_135_R[14]),
		.cost135_15(L_2_135_R[15]),
		.cost135_16(L_2_135_R[16]),
		.cost135_17(L_2_135_R[17]),
		.cost135_18(L_2_135_R[18]),
		.cost135_19(L_2_135_R[19]),
		.cost135_20(L_2_135_R[20]),
		.cost135_21(L_2_135_R[21]),
		.cost135_22(L_2_135_R[22]),
		.cost135_23(L_2_135_R[23]),
		.cost135_24(L_2_135_R[24]),
		.cost135_25(L_2_135_R[25]),
		.cost135_26(L_2_135_R[26]),
		.cost135_27(L_2_135_R[27]),
		.cost135_28(L_2_135_R[28]),
		.cost135_29(L_2_135_R[29]),
		.cost135_30(L_2_135_R[30]),
		.cost135_31(L_2_135_R[31]),
		.cost135_32(L_2_135_R[32]),
		.cost135_33(L_2_135_R[33]),
		.cost135_34(L_2_135_R[34]),
		.cost135_35(L_2_135_R[35]),
		.cost135_36(L_2_135_R[36]),
		.cost135_37(L_2_135_R[37]),
		.cost135_38(L_2_135_R[38]),
		.cost135_39(L_2_135_R[39]),
		.cost135_40(L_2_135_R[40]),
		.cost135_41(L_2_135_R[41]),
		.cost135_42(L_2_135_R[42]),
		.cost135_43(L_2_135_R[43]),
		.cost135_44(L_2_135_R[44]),
		.cost135_45(L_2_135_R[45]),
		.cost135_46(L_2_135_R[46]),
		.cost135_47(L_2_135_R[47]),
		.cost135_48(L_2_135_R[48]),
		.cost135_49(L_2_135_R[49]),
		.cost135_50(L_2_135_R[50]),
		.cost135_51(L_2_135_R[51]),
		.cost135_52(L_2_135_R[52]),
		.cost135_53(L_2_135_R[53]),
		.cost135_54(L_2_135_R[54]),
		.cost135_55(L_2_135_R[55]),
		.cost135_56(L_2_135_R[56]),
		.cost135_57(L_2_135_R[57]),
		.cost135_58(L_2_135_R[58]),
		.cost135_59(L_2_135_R[59]),
		.cost135_60(L_2_135_R[60]),
		.cost135_61(L_2_135_R[61]),
		.cost135_62(L_2_135_R[62]),
		.cost135_63(L_2_135_R[63]),
	
		.agg3_0_0(new3_L0_R[0]),
		.agg3_0_1(new3_L0_R[1]),
		.agg3_0_2(new3_L0_R[2]),
		.agg3_0_3(new3_L0_R[3]),
		.agg3_0_4(new3_L0_R[4]),
		.agg3_0_5(new3_L0_R[5]),
		.agg3_0_6(new3_L0_R[6]),
		.agg3_0_7(new3_L0_R[7]),
		.agg3_0_8(new3_L0_R[8]),
		.agg3_0_9(new3_L0_R[9]),
		.agg3_0_10(new3_L0_R[10]),
		.agg3_0_11(new3_L0_R[11]),
		.agg3_0_12(new3_L0_R[12]),
		.agg3_0_13(new3_L0_R[13]),
		.agg3_0_14(new3_L0_R[14]),
		.agg3_0_15(new3_L0_R[15]),
		.agg3_0_16(new3_L0_R[16]),
		.agg3_0_17(new3_L0_R[17]),
		.agg3_0_18(new3_L0_R[18]),
		.agg3_0_19(new3_L0_R[19]),
		.agg3_0_20(new3_L0_R[20]),
		.agg3_0_21(new3_L0_R[21]),
		.agg3_0_22(new3_L0_R[22]),
		.agg3_0_23(new3_L0_R[23]),
		.agg3_0_24(new3_L0_R[24]),
		.agg3_0_25(new3_L0_R[25]),
		.agg3_0_26(new3_L0_R[26]),
		.agg3_0_27(new3_L0_R[27]),
		.agg3_0_28(new3_L0_R[28]),
		.agg3_0_29(new3_L0_R[29]),
		.agg3_0_30(new3_L0_R[30]),
		.agg3_0_31(new3_L0_R[31]),
		.agg3_0_32(new3_L0_R[32]),
		.agg3_0_33(new3_L0_R[33]),
		.agg3_0_34(new3_L0_R[34]),
		.agg3_0_35(new3_L0_R[35]),
		.agg3_0_36(new3_L0_R[36]),
		.agg3_0_37(new3_L0_R[37]),
		.agg3_0_38(new3_L0_R[38]),
		.agg3_0_39(new3_L0_R[39]),
		.agg3_0_40(new3_L0_R[40]),
		.agg3_0_41(new3_L0_R[41]),
		.agg3_0_42(new3_L0_R[42]),
		.agg3_0_43(new3_L0_R[43]),
		.agg3_0_44(new3_L0_R[44]),
		.agg3_0_45(new3_L0_R[45]),
		.agg3_0_46(new3_L0_R[46]),
		.agg3_0_47(new3_L0_R[47]),
		.agg3_0_48(new3_L0_R[48]),
		.agg3_0_49(new3_L0_R[49]),
		.agg3_0_50(new3_L0_R[50]),
		.agg3_0_51(new3_L0_R[51]),
		.agg3_0_52(new3_L0_R[52]),
		.agg3_0_53(new3_L0_R[53]),
		.agg3_0_54(new3_L0_R[54]),
		.agg3_0_55(new3_L0_R[55]),
		.agg3_0_56(new3_L0_R[56]),
		.agg3_0_57(new3_L0_R[57]),
		.agg3_0_58(new3_L0_R[58]),
		.agg3_0_59(new3_L0_R[59]),
		.agg3_0_60(new3_L0_R[60]),
		.agg3_0_61(new3_L0_R[61]),
		.agg3_0_62(new3_L0_R[62]),
		.agg3_0_63(new3_L0_R[63]),
		
		.agg3_135_0(new3_L135_R[0]),
		.agg3_135_1(new3_L135_R[1]),
		.agg3_135_2(new3_L135_R[2]),
		.agg3_135_3(new3_L135_R[3]),
		.agg3_135_4(new3_L135_R[4]),
		.agg3_135_5(new3_L135_R[5]),
		.agg3_135_6(new3_L135_R[6]),
		.agg3_135_7(new3_L135_R[7]),
		.agg3_135_8(new3_L135_R[8]),
		.agg3_135_9(new3_L135_R[9]),
		.agg3_135_10(new3_L135_R[10]),
		.agg3_135_11(new3_L135_R[11]),
		.agg3_135_12(new3_L135_R[12]),
		.agg3_135_13(new3_L135_R[13]),
		.agg3_135_14(new3_L135_R[14]),
		.agg3_135_15(new3_L135_R[15]),
		.agg3_135_16(new3_L135_R[16]),
		.agg3_135_17(new3_L135_R[17]),
		.agg3_135_18(new3_L135_R[18]),
		.agg3_135_19(new3_L135_R[19]),
		.agg3_135_20(new3_L135_R[20]),
		.agg3_135_21(new3_L135_R[21]),
		.agg3_135_22(new3_L135_R[22]),
		.agg3_135_23(new3_L135_R[23]),
		.agg3_135_24(new3_L135_R[24]),
		.agg3_135_25(new3_L135_R[25]),
		.agg3_135_26(new3_L135_R[26]),
		.agg3_135_27(new3_L135_R[27]),
		.agg3_135_28(new3_L135_R[28]),
		.agg3_135_29(new3_L135_R[29]),
		.agg3_135_30(new3_L135_R[30]),
		.agg3_135_31(new3_L135_R[31]),
		.agg3_135_32(new3_L135_R[32]),
		.agg3_135_33(new3_L135_R[33]),
		.agg3_135_34(new3_L135_R[34]),
		.agg3_135_35(new3_L135_R[35]),
		.agg3_135_36(new3_L135_R[36]),
		.agg3_135_37(new3_L135_R[37]),
		.agg3_135_38(new3_L135_R[38]),
		.agg3_135_39(new3_L135_R[39]),
		.agg3_135_40(new3_L135_R[40]),
		.agg3_135_41(new3_L135_R[41]),
		.agg3_135_42(new3_L135_R[42]),
		.agg3_135_43(new3_L135_R[43]),
		.agg3_135_44(new3_L135_R[44]),
		.agg3_135_45(new3_L135_R[45]),
		.agg3_135_46(new3_L135_R[46]),
		.agg3_135_47(new3_L135_R[47]),
		.agg3_135_48(new3_L135_R[48]),
		.agg3_135_49(new3_L135_R[49]),
		.agg3_135_50(new3_L135_R[50]),
		.agg3_135_51(new3_L135_R[51]),
		.agg3_135_52(new3_L135_R[52]),
		.agg3_135_53(new3_L135_R[53]),
		.agg3_135_54(new3_L135_R[54]),
		.agg3_135_55(new3_L135_R[55]),
		.agg3_135_56(new3_L135_R[56]),
		.agg3_135_57(new3_L135_R[57]),
		.agg3_135_58(new3_L135_R[58]),
		.agg3_135_59(new3_L135_R[59]),
		.agg3_135_60(new3_L135_R[60]),
		.agg3_135_61(new3_L135_R[61]),
		.agg3_135_62(new3_L135_R[62]),
		.agg3_135_63(new3_L135_R[63]),
	
		.L0_0(L_3_0_R[0]),
		.L0_1(L_3_0_R[1]),
		.L0_2(L_3_0_R[2]),
		.L0_3(L_3_0_R[3]),
		.L0_4(L_3_0_R[4]),
		.L0_5(L_3_0_R[5]),
		.L0_6(L_3_0_R[6]),
		.L0_7(L_3_0_R[7]),
		.L0_8(L_3_0_R[8]),
		.L0_9(L_3_0_R[9]),
		.L0_10(L_3_0_R[10]),
		.L0_11(L_3_0_R[11]),
		.L0_12(L_3_0_R[12]),
		.L0_13(L_3_0_R[13]),
		.L0_14(L_3_0_R[14]),
		.L0_15(L_3_0_R[15]),
		.L0_16(L_3_0_R[16]),
		.L0_17(L_3_0_R[17]),
		.L0_18(L_3_0_R[18]),
		.L0_19(L_3_0_R[19]),
		.L0_20(L_3_0_R[20]),
		.L0_21(L_3_0_R[21]),
		.L0_22(L_3_0_R[22]),
		.L0_23(L_3_0_R[23]),
		.L0_24(L_3_0_R[24]),
		.L0_25(L_3_0_R[25]),
		.L0_26(L_3_0_R[26]),
		.L0_27(L_3_0_R[27]),
		.L0_28(L_3_0_R[28]),
		.L0_29(L_3_0_R[29]),
		.L0_30(L_3_0_R[30]),
		.L0_31(L_3_0_R[31]),
		.L0_32(L_3_0_R[32]),
		.L0_33(L_3_0_R[33]),
		.L0_34(L_3_0_R[34]),
		.L0_35(L_3_0_R[35]),
		.L0_36(L_3_0_R[36]),
		.L0_37(L_3_0_R[37]),
		.L0_38(L_3_0_R[38]),
		.L0_39(L_3_0_R[39]),
		.L0_40(L_3_0_R[40]),
		.L0_41(L_3_0_R[41]),
		.L0_42(L_3_0_R[42]),
		.L0_43(L_3_0_R[43]),
		.L0_44(L_3_0_R[44]),
		.L0_45(L_3_0_R[45]),
		.L0_46(L_3_0_R[46]),
		.L0_47(L_3_0_R[47]),
		.L0_48(L_3_0_R[48]),
		.L0_49(L_3_0_R[49]),
		.L0_50(L_3_0_R[50]),
		.L0_51(L_3_0_R[51]),
		.L0_52(L_3_0_R[52]),
		.L0_53(L_3_0_R[53]),
		.L0_54(L_3_0_R[54]),
		.L0_55(L_3_0_R[55]),
		.L0_56(L_3_0_R[56]),
		.L0_57(L_3_0_R[57]),
		.L0_58(L_3_0_R[58]),
		.L0_59(L_3_0_R[59]),
		.L0_60(L_3_0_R[60]),
		.L0_61(L_3_0_R[61]),
		.L0_62(L_3_0_R[62]),
		.L0_63(L_3_0_R[63]),
	
		.L135_0(L_3_135_R[0]),
		.L135_1(L_3_135_R[1]),
		.L135_2(L_3_135_R[2]),
		.L135_3(L_3_135_R[3]),
		.L135_4(L_3_135_R[4]),
		.L135_5(L_3_135_R[5]),
		.L135_6(L_3_135_R[6]),
		.L135_7(L_3_135_R[7]),
		.L135_8(L_3_135_R[8]),
		.L135_9(L_3_135_R[9]),
		.L135_10(L_3_135_R[10]),
		.L135_11(L_3_135_R[11]),
		.L135_12(L_3_135_R[12]),
		.L135_13(L_3_135_R[13]),
		.L135_14(L_3_135_R[14]),
		.L135_15(L_3_135_R[15]),
		.L135_16(L_3_135_R[16]),
		.L135_17(L_3_135_R[17]),
		.L135_18(L_3_135_R[18]),
		.L135_19(L_3_135_R[19]),
		.L135_20(L_3_135_R[20]),
		.L135_21(L_3_135_R[21]),
		.L135_22(L_3_135_R[22]),
		.L135_23(L_3_135_R[23]),
		.L135_24(L_3_135_R[24]),
		.L135_25(L_3_135_R[25]),
		.L135_26(L_3_135_R[26]),
		.L135_27(L_3_135_R[27]),
		.L135_28(L_3_135_R[28]),
		.L135_29(L_3_135_R[29]),
		.L135_30(L_3_135_R[30]),
		.L135_31(L_3_135_R[31]),
		.L135_32(L_3_135_R[32]),
		.L135_33(L_3_135_R[33]),
		.L135_34(L_3_135_R[34]),
		.L135_35(L_3_135_R[35]),
		.L135_36(L_3_135_R[36]),
		.L135_37(L_3_135_R[37]),
		.L135_38(L_3_135_R[38]),
		.L135_39(L_3_135_R[39]),
		.L135_40(L_3_135_R[40]),
		.L135_41(L_3_135_R[41]),
		.L135_42(L_3_135_R[42]),
		.L135_43(L_3_135_R[43]),
		.L135_44(L_3_135_R[44]),
		.L135_45(L_3_135_R[45]),
		.L135_46(L_3_135_R[46]),
		.L135_47(L_3_135_R[47]),
		.L135_48(L_3_135_R[48]),
		.L135_49(L_3_135_R[49]),
		.L135_50(L_3_135_R[50]),
		.L135_51(L_3_135_R[51]),
		.L135_52(L_3_135_R[52]),
		.L135_53(L_3_135_R[53]),
		.L135_54(L_3_135_R[54]),
		.L135_55(L_3_135_R[55]),
		.L135_56(L_3_135_R[56]),
		.L135_57(L_3_135_R[57]),
		.L135_58(L_3_135_R[58]),
		.L135_59(L_3_135_R[59]),
		.L135_60(L_3_135_R[60]),
		.L135_61(L_3_135_R[61]),
		.L135_62(L_3_135_R[62]),
		.L135_63(L_3_135_R[63])    
		);
	
	//0
	
	wire [(cost_width*8-1):0] din_0_R_1 = {L_0_R[7][0],L_0_R[6][0],L_0_R[5][0],L_0_R[4][0],L_0_R[3][0],L_0_R[2][0],L_0_R[1][0],L_0_R[0][0]};
	wire [(cost_width*8-1):0] din_0_R_2 = {L_0_R[15][0],L_0_R[14][0],L_0_R[13][0],L_0_R[12][0],L_0_R[11][0],L_0_R[10][0],L_0_R[9][0],L_0_R[8][0]};
	wire [(cost_width*8-1):0] din_0_R_3 = {L_0_R[23][0],L_0_R[22][0],L_0_R[21][0],L_0_R[20][0],L_0_R[19][0],L_0_R[18][0],L_0_R[17][0],L_0_R[16][0]};
	wire [(cost_width*8-1):0] din_0_R_4 = {L_0_R[31][0],L_0_R[30][0],L_0_R[29][0],L_0_R[28][0],L_0_R[27][0],L_0_R[26][0],L_0_R[25][0],L_0_R[24][0]};
	wire [(cost_width*8-1):0] din_0_R_5 = {L_0_R[39][0],L_0_R[38][0],L_0_R[37][0],L_0_R[36][0],L_0_R[35][0],L_0_R[34][0],L_0_R[33][0],L_0_R[32][0]};
	wire [(cost_width*8-1):0] din_0_R_6 = {L_0_R[47][0],L_0_R[46][0],L_0_R[45][0],L_0_R[44][0],L_0_R[43][0],L_0_R[42][0],L_0_R[41][0],L_0_R[40][0]};
	wire [(cost_width*8-1):0] din_0_R_7 = {L_0_R[55][0],L_0_R[54][0],L_0_R[53][0],L_0_R[52][0],L_0_R[51][0],L_0_R[50][0],L_0_R[49][0],L_0_R[48][0]};
	wire [(cost_width*8-1):0] din_0_R_8 = {L_0_R[63][0],L_0_R[62][0],L_0_R[61][0],L_0_R[60][0],L_0_R[59][0],L_0_R[58][0],L_0_R[57][0],L_0_R[56][0]};
	
	wire [(cost_width*64-1):0] din_0_R = {din_0_R_8,din_0_R_7,din_0_R_6,din_0_R_5,din_0_R_4,din_0_R_3,din_0_R_2,din_0_R_1};
	wire [(cost_width*64-1):0] dout_0_R = Q_Aggregation0_Ram_2[(cost_width*64-1):0];

	genvar i;
	generate for(i=0;i<64;i=i+1) begin: loop
			assign L_0_R[i][1] = dout_0_R[i*cost_width+(cost_width-1):i*cost_width];
		end
	endgenerate
	
	//135
	wire [((cost_width-2)*8-1):0] din_135_R_1 = {L_135_R[7][0],L_135_R[6][0],L_135_R[5][0],L_135_R[4][0],L_135_R[3][0],L_135_R[2][0],L_135_R[1][0],L_135_R[0][0]};
	wire [((cost_width-2)*8-1):0] din_135_R_2 = {L_135_R[15][0],L_135_R[14][0],L_135_R[13][0],L_135_R[12][0],L_135_R[11][0],L_135_R[10][0],L_135_R[9][0],L_135_R[8][0]};
	wire [((cost_width-2)*8-1):0] din_135_R_3 = {L_135_R[23][0],L_135_R[22][0],L_135_R[21][0],L_135_R[20][0],L_135_R[19][0],L_135_R[18][0],L_135_R[17][0],L_135_R[16][0]};
	wire [((cost_width-2)*8-1):0] din_135_R_4 = {L_135_R[31][0],L_135_R[30][0],L_135_R[29][0],L_135_R[28][0],L_135_R[27][0],L_135_R[26][0],L_135_R[25][0],L_135_R[24][0]};
	wire [((cost_width-2)*8-1):0] din_135_R_5 = {L_135_R[39][0],L_135_R[38][0],L_135_R[37][0],L_135_R[36][0],L_135_R[35][0],L_135_R[34][0],L_135_R[33][0],L_135_R[32][0]};
	wire [((cost_width-2)*8-1):0] din_135_R_6 = {L_135_R[47][0],L_135_R[46][0],L_135_R[45][0],L_135_R[44][0],L_135_R[43][0],L_135_R[42][0],L_135_R[41][0],L_135_R[40][0]};
	wire [((cost_width-2)*8-1):0] din_135_R_7 = {L_135_R[55][0],L_135_R[54][0],L_135_R[53][0],L_135_R[52][0],L_135_R[51][0],L_135_R[50][0],L_135_R[49][0],L_135_R[48][0]};
	wire [((cost_width-2)*8-1):0] din_135_R_8 = {L_135_R[63][0],L_135_R[62][0],L_135_R[61][0],L_135_R[60][0],L_135_R[59][0],L_135_R[58][0],L_135_R[57][0],L_135_R[56][0]};
	wire [((cost_width-2)*64-1):0]din_135_R = {din_135_R_8,din_135_R_7,din_135_R_6,din_135_R_5,din_135_R_4,din_135_R_3,din_135_R_2,din_135_R_1};
	wire [((cost_width-2)*64-1):0] dout_135_R = Q_Aggregation135_Ram_2[((cost_width-2)*64-1):0];

	genvar j;
	generate for(j=0;j<64;j=j+1) begin: loop2
			assign L_135_R[j][1] = dout_135_R[j*(cost_width-2)+(cost_width-3):j*(cost_width-2)];
		end
	endgenerate
	
	//Aggregation modules for the right direction		
	agg2#(cost_width) agg2_Right(
		.clk(clk),
		.rst(rst),
		.clken(clken0),
		.en_first(en_first_R_agg2),

        .P1({P1,2'b00}),
        .P2({P2,2'b00}),
		
		.agg0_0(L_0_R[0][2]),
		.agg0_1(L_0_R[1][2]),
		.agg0_2(L_0_R[2][2]),
		.agg0_3(L_0_R[3][2]),
		.agg0_4(L_0_R[4][2]),
		.agg0_5(L_0_R[5][2]),
		.agg0_6(L_0_R[6][2]),
		.agg0_7(L_0_R[7][2]),
		.agg0_8(L_0_R[8][2]),
		.agg0_9(L_0_R[9][2]),
		.agg0_10(L_0_R[10][2]),
		.agg0_11(L_0_R[11][2]),
		.agg0_12(L_0_R[12][2]),
		.agg0_13(L_0_R[13][2]),
		.agg0_14(L_0_R[14][2]),
		.agg0_15(L_0_R[15][2]),
		.agg0_16(L_0_R[16][2]),
		.agg0_17(L_0_R[17][2]),
		.agg0_18(L_0_R[18][2]),
		.agg0_19(L_0_R[19][2]),
		.agg0_20(L_0_R[20][2]),
		.agg0_21(L_0_R[21][2]),
		.agg0_22(L_0_R[22][2]),
		.agg0_23(L_0_R[23][2]),
		.agg0_24(L_0_R[24][2]),
		.agg0_25(L_0_R[25][2]),
		.agg0_26(L_0_R[26][2]),
		.agg0_27(L_0_R[27][2]),
		.agg0_28(L_0_R[28][2]),
		.agg0_29(L_0_R[29][2]),
		.agg0_30(L_0_R[30][2]),
		.agg0_31(L_0_R[31][2]),
		.agg0_32(L_0_R[32][2]),
		.agg0_33(L_0_R[33][2]),
		.agg0_34(L_0_R[34][2]),
		.agg0_35(L_0_R[35][2]),
		.agg0_36(L_0_R[36][2]),
		.agg0_37(L_0_R[37][2]),
		.agg0_38(L_0_R[38][2]),
		.agg0_39(L_0_R[39][2]),
		.agg0_40(L_0_R[40][2]),
		.agg0_41(L_0_R[41][2]),
		.agg0_42(L_0_R[42][2]),
		.agg0_43(L_0_R[43][2]),
		.agg0_44(L_0_R[44][2]),
		.agg0_45(L_0_R[45][2]),
		.agg0_46(L_0_R[46][2]),
		.agg0_47(L_0_R[47][2]),
		.agg0_48(L_0_R[48][2]),
		.agg0_49(L_0_R[49][2]),
		.agg0_50(L_0_R[50][2]),
		.agg0_51(L_0_R[51][2]),
		.agg0_52(L_0_R[52][2]),
		.agg0_53(L_0_R[53][2]),
		.agg0_54(L_0_R[54][2]),
		.agg0_55(L_0_R[55][2]),
		.agg0_56(L_0_R[56][2]),
		.agg0_57(L_0_R[57][2]),
		.agg0_58(L_0_R[58][2]),
		.agg0_59(L_0_R[59][2]),
		.agg0_60(L_0_R[60][2]),
		.agg0_61(L_0_R[61][2]),
		.agg0_62(L_0_R[62][2]),
		.agg0_63(L_0_R[63][2]),
	
		.cost0_0(L_0_R[0][1]),
		.cost0_1(L_0_R[1][1]),
		.cost0_2(L_0_R[2][1]),
		.cost0_3(L_0_R[3][1]),
		.cost0_4(L_0_R[4][1]),
		.cost0_5(L_0_R[5][1]),
		.cost0_6(L_0_R[6][1]),
		.cost0_7(L_0_R[7][1]),
		.cost0_8(L_0_R[8][1]),
		.cost0_9(L_0_R[9][1]),
		.cost0_10(L_0_R[10][1]),
		.cost0_11(L_0_R[11][1]),
		.cost0_12(L_0_R[12][1]),
		.cost0_13(L_0_R[13][1]),
		.cost0_14(L_0_R[14][1]),
		.cost0_15(L_0_R[15][1]),
		.cost0_16(L_0_R[16][1]),
		.cost0_17(L_0_R[17][1]),
		.cost0_18(L_0_R[18][1]),
		.cost0_19(L_0_R[19][1]),
		.cost0_20(L_0_R[20][1]),
		.cost0_21(L_0_R[21][1]),
		.cost0_22(L_0_R[22][1]),
		.cost0_23(L_0_R[23][1]),
		.cost0_24(L_0_R[24][1]),
		.cost0_25(L_0_R[25][1]),
		.cost0_26(L_0_R[26][1]),
		.cost0_27(L_0_R[27][1]),
		.cost0_28(L_0_R[28][1]),
		.cost0_29(L_0_R[29][1]),
		.cost0_30(L_0_R[30][1]),
		.cost0_31(L_0_R[31][1]),
		.cost0_32(L_0_R[32][1]),
		.cost0_33(L_0_R[33][1]),
		.cost0_34(L_0_R[34][1]),
		.cost0_35(L_0_R[35][1]),
		.cost0_36(L_0_R[36][1]),
		.cost0_37(L_0_R[37][1]),
		.cost0_38(L_0_R[38][1]),
		.cost0_39(L_0_R[39][1]),
		.cost0_40(L_0_R[40][1]),
		.cost0_41(L_0_R[41][1]),
		.cost0_42(L_0_R[42][1]),
		.cost0_43(L_0_R[43][1]),
		.cost0_44(L_0_R[44][1]),
		.cost0_45(L_0_R[45][1]),
		.cost0_46(L_0_R[46][1]),
		.cost0_47(L_0_R[47][1]),
		.cost0_48(L_0_R[48][1]),
		.cost0_49(L_0_R[49][1]),
		.cost0_50(L_0_R[50][1]),
		.cost0_51(L_0_R[51][1]),
		.cost0_52(L_0_R[52][1]),
		.cost0_53(L_0_R[53][1]),
		.cost0_54(L_0_R[54][1]),
		.cost0_55(L_0_R[55][1]),
		.cost0_56(L_0_R[56][1]),
		.cost0_57(L_0_R[57][1]),
		.cost0_58(L_0_R[58][1]),
		.cost0_59(L_0_R[59][1]),
		.cost0_60(L_0_R[60][1]),
		.cost0_61(L_0_R[61][1]),
		.cost0_62(L_0_R[62][1]),
		.cost0_63(L_0_R[63][1]),
	
		.cost135_0(L_135_R[0][1]),
		.cost135_1(L_135_R[1][1]),
		.cost135_2(L_135_R[2][1]),
		.cost135_3(L_135_R[3][1]),
		.cost135_4(L_135_R[4][1]),
		.cost135_5(L_135_R[5][1]),
		.cost135_6(L_135_R[6][1]),
		.cost135_7(L_135_R[7][1]),
		.cost135_8(L_135_R[8][1]),
		.cost135_9(L_135_R[9][1]),
		.cost135_10(L_135_R[10][1]),
		.cost135_11(L_135_R[11][1]),
		.cost135_12(L_135_R[12][1]),
		.cost135_13(L_135_R[13][1]),
		.cost135_14(L_135_R[14][1]),
		.cost135_15(L_135_R[15][1]),
		.cost135_16(L_135_R[16][1]),
		.cost135_17(L_135_R[17][1]),
		.cost135_18(L_135_R[18][1]),
		.cost135_19(L_135_R[19][1]),
		.cost135_20(L_135_R[20][1]),
		.cost135_21(L_135_R[21][1]),
		.cost135_22(L_135_R[22][1]),
		.cost135_23(L_135_R[23][1]),
		.cost135_24(L_135_R[24][1]),
		.cost135_25(L_135_R[25][1]),
		.cost135_26(L_135_R[26][1]),
		.cost135_27(L_135_R[27][1]),	
		.cost135_28(L_135_R[28][1]),
		.cost135_29(L_135_R[29][1]),
		.cost135_30(L_135_R[30][1]),
		.cost135_31(L_135_R[31][1]),	
		.cost135_32(L_135_R[32][1]),
		.cost135_33(L_135_R[33][1]),
		.cost135_34(L_135_R[34][1]),
		.cost135_35(L_135_R[35][1]),
		.cost135_36(L_135_R[36][1]),
		.cost135_37(L_135_R[37][1]),
		.cost135_38(L_135_R[38][1]),
		.cost135_39(L_135_R[39][1]),
		.cost135_40(L_135_R[40][1]),
		.cost135_41(L_135_R[41][1]),
		.cost135_42(L_135_R[42][1]),
		.cost135_43(L_135_R[43][1]),
		.cost135_44(L_135_R[44][1]),
		.cost135_45(L_135_R[45][1]),
		.cost135_46(L_135_R[46][1]),
		.cost135_47(L_135_R[47][1]),
		.cost135_48(L_135_R[48][1]),
		.cost135_49(L_135_R[49][1]),
		.cost135_50(L_135_R[50][1]),
		.cost135_51(L_135_R[51][1]),
		.cost135_52(L_135_R[52][1]),
		.cost135_53(L_135_R[53][1]),
		.cost135_54(L_135_R[54][1]),
		.cost135_55(L_135_R[55][1]),
		.cost135_56(L_135_R[56][1]),
		.cost135_57(L_135_R[57][1]),	
		.cost135_58(L_135_R[58][1]),
		.cost135_59(L_135_R[59][1]),
		.cost135_60(L_135_R[60][1]),
		.cost135_61(L_135_R[61][1]),
		.cost135_62(L_135_R[62][1]),
		.cost135_63(L_135_R[63][1]),
	
		.min_0_in(min_0_R),
		.min_135(min_135_R),
		.min_0_out(min_0_R),
	
		.L0_0(L_0_R[0][2]),
		.L0_1(L_0_R[1][2]),
		.L0_2(L_0_R[2][2]),
		.L0_3(L_0_R[3][2]),
		.L0_4(L_0_R[4][2]),
		.L0_5(L_0_R[5][2]),
		.L0_6(L_0_R[6][2]),
		.L0_7(L_0_R[7][2]),
		.L0_8(L_0_R[8][2]),
		.L0_9(L_0_R[9][2]),
		.L0_10(L_0_R[10][2]),
		.L0_11(L_0_R[11][2]),
		.L0_12(L_0_R[12][2]),
		.L0_13(L_0_R[13][2]),
		.L0_14(L_0_R[14][2]),
		.L0_15(L_0_R[15][2]),
		.L0_16(L_0_R[16][2]),
		.L0_17(L_0_R[17][2]),
		.L0_18(L_0_R[18][2]),
		.L0_19(L_0_R[19][2]),
		.L0_20(L_0_R[20][2]),
		.L0_21(L_0_R[21][2]),
		.L0_22(L_0_R[22][2]),
		.L0_23(L_0_R[23][2]),
		.L0_24(L_0_R[24][2]),
		.L0_25(L_0_R[25][2]),
		.L0_26(L_0_R[26][2]),
		.L0_27(L_0_R[27][2]),
		.L0_28(L_0_R[28][2]),
		.L0_29(L_0_R[29][2]),
		.L0_30(L_0_R[30][2]),
		.L0_31(L_0_R[31][2]),
		.L0_32(L_0_R[32][2]),
		.L0_33(L_0_R[33][2]),
		.L0_34(L_0_R[34][2]),
		.L0_35(L_0_R[35][2]),
		.L0_36(L_0_R[36][2]),
		.L0_37(L_0_R[37][2]),
		.L0_38(L_0_R[38][2]),
		.L0_39(L_0_R[39][2]),
		.L0_40(L_0_R[40][2]),
		.L0_41(L_0_R[41][2]),
		.L0_42(L_0_R[42][2]),
		.L0_43(L_0_R[43][2]),
		.L0_44(L_0_R[44][2]),
		.L0_45(L_0_R[45][2]),
		.L0_46(L_0_R[46][2]),
		.L0_47(L_0_R[47][2]),
		.L0_48(L_0_R[48][2]),
		.L0_49(L_0_R[49][2]),
		.L0_50(L_0_R[50][2]),
		.L0_51(L_0_R[51][2]),
		.L0_52(L_0_R[52][2]),
		.L0_53(L_0_R[53][2]),
		.L0_54(L_0_R[54][2]),
		.L0_55(L_0_R[55][2]),
		.L0_56(L_0_R[56][2]),
		.L0_57(L_0_R[57][2]),
		.L0_58(L_0_R[58][2]),
		.L0_59(L_0_R[59][2]),
		.L0_60(L_0_R[60][2]),
		.L0_61(L_0_R[61][2]),
		.L0_62(L_0_R[62][2]),
		.L0_63(L_0_R[63][2]),
	
		.L135_0(L_135_R[0][2]),
		.L135_1(L_135_R[1][2]),
		.L135_2(L_135_R[2][2]),
		.L135_3(L_135_R[3][2]),
		.L135_4(L_135_R[4][2]),
		.L135_5(L_135_R[5][2]),
		.L135_6(L_135_R[6][2]),
		.L135_7(L_135_R[7][2]),
		.L135_8(L_135_R[8][2]),
		.L135_9(L_135_R[9][2]),
		.L135_10(L_135_R[10][2]),
		.L135_11(L_135_R[11][2]),
		.L135_12(L_135_R[12][2]),
		.L135_13(L_135_R[13][2]),
		.L135_14(L_135_R[14][2]),
		.L135_15(L_135_R[15][2]),
		.L135_16(L_135_R[16][2]),
		.L135_17(L_135_R[17][2]),
		.L135_18(L_135_R[18][2]),
		.L135_19(L_135_R[19][2]),
		.L135_20(L_135_R[20][2]),
		.L135_21(L_135_R[21][2]),
		.L135_22(L_135_R[22][2]),
		.L135_23(L_135_R[23][2]),
		.L135_24(L_135_R[24][2]),
		.L135_25(L_135_R[25][2]),
		.L135_26(L_135_R[26][2]),
		.L135_27(L_135_R[27][2]),	
		.L135_28(L_135_R[28][2]),
		.L135_29(L_135_R[29][2]),
		.L135_30(L_135_R[30][2]),
		.L135_31(L_135_R[31][2]),
		.L135_32(L_135_R[32][2]),
		.L135_33(L_135_R[33][2]),
		.L135_34(L_135_R[34][2]),
		.L135_35(L_135_R[35][2]),
		.L135_36(L_135_R[36][2]),
		.L135_37(L_135_R[37][2]),
		.L135_38(L_135_R[38][2]),
		.L135_39(L_135_R[39][2]),
		.L135_40(L_135_R[40][2]),
		.L135_41(L_135_R[41][2]),
		.L135_42(L_135_R[42][2]),
		.L135_43(L_135_R[43][2]),
		.L135_44(L_135_R[44][2]),
		.L135_45(L_135_R[45][2]),
		.L135_46(L_135_R[46][2]),
		.L135_47(L_135_R[47][2]),
		.L135_48(L_135_R[48][2]),
		.L135_49(L_135_R[49][2]),
		.L135_50(L_135_R[50][2]),
		.L135_51(L_135_R[51][2]),
		.L135_52(L_135_R[52][2]),
		.L135_53(L_135_R[53][2]),
		.L135_54(L_135_R[54][2]),
		.L135_55(L_135_R[55][2]),
		.L135_56(L_135_R[56][2]),
		.L135_57(L_135_R[57][2]),	
		.L135_58(L_135_R[58][2]),
		.L135_59(L_135_R[59][2]),
		.L135_60(L_135_R[60][2]),
		.L135_61(L_135_R[61][2]),
		.L135_62(L_135_R[62][2]),
		.L135_63(L_135_R[63][2]),
		
		.cost_valid(cost_valid)
		);
	
	agg4#(cost_width) agg4_Right(
		.clk(clk),
		.rst0(rst0_R),
		.rst(rst),
		.clken(clken0),
		.en_first(en_first_R),//first pixel of every row
		.en_agg4(en_agg4_R),  //when second row comes
		.L0_0(cost_R_in[0]),
		.L0_1(cost_R_in[1]),
		.L0_2(cost_R_in[2]),
		.L0_3(cost_R_in[3]),
		.L0_4(cost_R_in[4]),
		.L0_5(cost_R_in[5]),
		.L0_6(cost_R_in[6]),
		.L0_7(cost_R_in[7]),
		.L0_8(cost_R_in[8]),
		.L0_9(cost_R_in[9]),
		.L0_10(cost_R_in[10]),
		.L0_11(cost_R_in[11]),
		.L0_12(cost_R_in[12]),
		.L0_13(cost_R_in[13]),
		.L0_14(cost_R_in[14]),
		.L0_15(cost_R_in[15]),
		.L0_16(cost_R_in[16]),
		.L0_17(cost_R_in[17]),
		.L0_18(cost_R_in[18]),
		.L0_19(cost_R_in[19]),
		.L0_20(cost_R_in[20]),
		.L0_21(cost_R_in[21]),
		.L0_22(cost_R_in[22]),
		.L0_23(cost_R_in[23]),
		.L0_24(cost_R_in[24]),
		.L0_25(cost_R_in[25]),
		.L0_26(cost_R_in[26]),
		.L0_27(cost_R_in[27]),
		.L0_28(cost_R_in[28]),
		.L0_29(cost_R_in[29]),
		.L0_30(cost_R_in[30]),
		.L0_31(cost_R_in[31]),
		.L0_32(cost_R_in[32]),
		.L0_33(cost_R_in[33]),
		.L0_34(cost_R_in[34]),
		.L0_35(cost_R_in[35]),
		.L0_36(cost_R_in[36]),
		.L0_37(cost_R_in[37]),
		.L0_38(cost_R_in[38]),
		.L0_39(cost_R_in[39]),
		.L0_40(cost_R_in[40]),
		.L0_41(cost_R_in[41]),
		.L0_42(cost_R_in[42]),
		.L0_43(cost_R_in[43]),
		.L0_44(cost_R_in[44]),
		.L0_45(cost_R_in[45]),
		.L0_46(cost_R_in[46]),
		.L0_47(cost_R_in[47]),
		.L0_48(cost_R_in[48]),
		.L0_49(cost_R_in[49]),
		.L0_50(cost_R_in[50]),
		.L0_51(cost_R_in[51]),
		.L0_52(cost_R_in[52]),
		.L0_53(cost_R_in[53]),
		.L0_54(cost_R_in[54]),
		.L0_55(cost_R_in[55]),
		.L0_56(cost_R_in[56]),
		.L0_57(cost_R_in[57]),
		.L0_58(cost_R_in[58]),
		.L0_59(cost_R_in[59]),
		.L0_60(cost_R_in[60]),
		.L0_61(cost_R_in[61]),
		.L0_62(cost_R_in[62]),
		.L0_63(cost_R_in[63]),
	
		.L135_0(cost_R_in[0][cost_width-1:2]),
		.L135_1(cost_R_in[1][cost_width-1:2]),
		.L135_2(cost_R_in[2][cost_width-1:2]),
		.L135_3(cost_R_in[3][cost_width-1:2]),
		.L135_4(cost_R_in[4][cost_width-1:2]),
		.L135_5(cost_R_in[5][cost_width-1:2]),
		.L135_6(cost_R_in[6][cost_width-1:2]),
		.L135_7(cost_R_in[7][cost_width-1:2]),
		.L135_8(cost_R_in[8][cost_width-1:2]),
		.L135_9(cost_R_in[9][cost_width-1:2]),
		.L135_10(cost_R_in[10][cost_width-1:2]),
		.L135_11(cost_R_in[11][cost_width-1:2]),
		.L135_12(cost_R_in[12][cost_width-1:2]),
		.L135_13(cost_R_in[13][cost_width-1:2]),
		.L135_14(cost_R_in[14][cost_width-1:2]),
		.L135_15(cost_R_in[15][cost_width-1:2]),
		.L135_16(cost_R_in[16][cost_width-1:2]),
		.L135_17(cost_R_in[17][cost_width-1:2]),
		.L135_18(cost_R_in[18][cost_width-1:2]),
		.L135_19(cost_R_in[19][cost_width-1:2]),
		.L135_20(cost_R_in[20][cost_width-1:2]),
		.L135_21(cost_R_in[21][cost_width-1:2]),
		.L135_22(cost_R_in[22][cost_width-1:2]),
		.L135_23(cost_R_in[23][cost_width-1:2]),
		.L135_24(cost_R_in[24][cost_width-1:2]),
		.L135_25(cost_R_in[25][cost_width-1:2]),
		.L135_26(cost_R_in[26][cost_width-1:2]),
		.L135_27(cost_R_in[27][cost_width-1:2]),
		.L135_28(cost_R_in[28][cost_width-1:2]),
		.L135_29(cost_R_in[29][cost_width-1:2]),
		.L135_30(cost_R_in[30][cost_width-1:2]),
		.L135_31(cost_R_in[31][cost_width-1:2]),
		.L135_32(cost_R_in[32][cost_width-1:2]),
		.L135_33(cost_R_in[33][cost_width-1:2]),
		.L135_34(cost_R_in[34][cost_width-1:2]),
		.L135_35(cost_R_in[35][cost_width-1:2]),
		.L135_36(cost_R_in[36][cost_width-1:2]),
		.L135_37(cost_R_in[37][cost_width-1:2]),
		.L135_38(cost_R_in[38][cost_width-1:2]),
		.L135_39(cost_R_in[39][cost_width-1:2]),
		.L135_40(cost_R_in[40][cost_width-1:2]),
		.L135_41(cost_R_in[41][cost_width-1:2]),
		.L135_42(cost_R_in[42][cost_width-1:2]),
		.L135_43(cost_R_in[43][cost_width-1:2]),
		.L135_44(cost_R_in[44][cost_width-1:2]),
		.L135_45(cost_R_in[45][cost_width-1:2]),
		.L135_46(cost_R_in[46][cost_width-1:2]),
		.L135_47(cost_R_in[47][cost_width-1:2]),
		.L135_48(cost_R_in[48][cost_width-1:2]),
		.L135_49(cost_R_in[49][cost_width-1:2]),
		.L135_50(cost_R_in[50][cost_width-1:2]),
		.L135_51(cost_R_in[51][cost_width-1:2]),
		.L135_52(cost_R_in[52][cost_width-1:2]),
		.L135_53(cost_R_in[53][cost_width-1:2]),
		.L135_54(cost_R_in[54][cost_width-1:2]),
		.L135_55(cost_R_in[55][cost_width-1:2]),
		.L135_56(cost_R_in[56][cost_width-1:2]),
		.L135_57(cost_R_in[57][cost_width-1:2]),
		.L135_58(cost_R_in[58][cost_width-1:2]),
		.L135_59(cost_R_in[59][cost_width-1:2]),
		.L135_60(cost_R_in[60][cost_width-1:2]),
		.L135_61(cost_R_in[61][cost_width-1:2]),
		.L135_62(cost_R_in[62][cost_width-1:2]),
		.L135_63(cost_R_in[63][cost_width-1:2]),
	
		.new_L0_0(new4_L0_R[0]),
		.new_L0_1(new4_L0_R[1]),
		.new_L0_2(new4_L0_R[2]),
		.new_L0_3(new4_L0_R[3]),
		.new_L0_4(new4_L0_R[4]),
		.new_L0_5(new4_L0_R[5]),
		.new_L0_6(new4_L0_R[6]),
		.new_L0_7(new4_L0_R[7]),
		.new_L0_8(new4_L0_R[8]),
		.new_L0_9(new4_L0_R[9]),
		.new_L0_10(new4_L0_R[10]),
		.new_L0_11(new4_L0_R[11]),
		.new_L0_12(new4_L0_R[12]),
		.new_L0_13(new4_L0_R[13]),
		.new_L0_14(new4_L0_R[14]),
		.new_L0_15(new4_L0_R[15]),
		.new_L0_16(new4_L0_R[16]),
		.new_L0_17(new4_L0_R[17]),
		.new_L0_18(new4_L0_R[18]),
		.new_L0_19(new4_L0_R[19]),
		.new_L0_20(new4_L0_R[20]),
		.new_L0_21(new4_L0_R[21]),
		.new_L0_22(new4_L0_R[22]),
		.new_L0_23(new4_L0_R[23]),
		.new_L0_24(new4_L0_R[24]),
		.new_L0_25(new4_L0_R[25]),
		.new_L0_26(new4_L0_R[26]),
		.new_L0_27(new4_L0_R[27]),
		.new_L0_28(new4_L0_R[28]),
		.new_L0_29(new4_L0_R[29]),
		.new_L0_30(new4_L0_R[30]),
		.new_L0_31(new4_L0_R[31]),
		.new_L0_32(new4_L0_R[32]),
		.new_L0_33(new4_L0_R[33]),
		.new_L0_34(new4_L0_R[34]),
		.new_L0_35(new4_L0_R[35]),
		.new_L0_36(new4_L0_R[36]),
		.new_L0_37(new4_L0_R[37]),
		.new_L0_38(new4_L0_R[38]),
		.new_L0_39(new4_L0_R[39]),
		.new_L0_40(new4_L0_R[40]),
		.new_L0_41(new4_L0_R[41]),
		.new_L0_42(new4_L0_R[42]),
		.new_L0_43(new4_L0_R[43]),
		.new_L0_44(new4_L0_R[44]),
		.new_L0_45(new4_L0_R[45]),
		.new_L0_46(new4_L0_R[46]),
		.new_L0_47(new4_L0_R[47]),
		.new_L0_48(new4_L0_R[48]),
		.new_L0_49(new4_L0_R[49]),
		.new_L0_50(new4_L0_R[50]),
		.new_L0_51(new4_L0_R[51]),
		.new_L0_52(new4_L0_R[52]),
		.new_L0_53(new4_L0_R[53]),
		.new_L0_54(new4_L0_R[54]),
		.new_L0_55(new4_L0_R[55]),
		.new_L0_56(new4_L0_R[56]),
		.new_L0_57(new4_L0_R[57]),
		.new_L0_58(new4_L0_R[58]),
		.new_L0_59(new4_L0_R[59]),
		.new_L0_60(new4_L0_R[60]),
		.new_L0_61(new4_L0_R[61]),
		.new_L0_62(new4_L0_R[62]),
		.new_L0_63(new4_L0_R[63]),	
		
		.new_L135_0(new4_L135_R[0]),
		.new_L135_1(new4_L135_R[1]),
		.new_L135_2(new4_L135_R[2]),
		.new_L135_3(new4_L135_R[3]),
		.new_L135_4(new4_L135_R[4]),
		.new_L135_5(new4_L135_R[5]),
		.new_L135_6(new4_L135_R[6]),
		.new_L135_7(new4_L135_R[7]),
		.new_L135_8(new4_L135_R[8]),
		.new_L135_9(new4_L135_R[9]),
		.new_L135_10(new4_L135_R[10]),
		.new_L135_11(new4_L135_R[11]),
		.new_L135_12(new4_L135_R[12]),
		.new_L135_13(new4_L135_R[13]),
		.new_L135_14(new4_L135_R[14]),
		.new_L135_15(new4_L135_R[15]),
		.new_L135_16(new4_L135_R[16]),
		.new_L135_17(new4_L135_R[17]),
		.new_L135_18(new4_L135_R[18]),
		.new_L135_19(new4_L135_R[19]),
		.new_L135_20(new4_L135_R[20]),
		.new_L135_21(new4_L135_R[21]),
		.new_L135_22(new4_L135_R[22]),
		.new_L135_23(new4_L135_R[23]),
		.new_L135_24(new4_L135_R[24]),
		.new_L135_25(new4_L135_R[25]),
		.new_L135_26(new4_L135_R[26]),
		.new_L135_27(new4_L135_R[27]),
		.new_L135_28(new4_L135_R[28]),
		.new_L135_29(new4_L135_R[29]),
		.new_L135_30(new4_L135_R[30]),
		.new_L135_31(new4_L135_R[31]),
		.new_L135_32(new4_L135_R[32]),
		.new_L135_33(new4_L135_R[33]),
		.new_L135_34(new4_L135_R[34]),
		.new_L135_35(new4_L135_R[35]),
		.new_L135_36(new4_L135_R[36]),
		.new_L135_37(new4_L135_R[37]),
		.new_L135_38(new4_L135_R[38]),
		.new_L135_39(new4_L135_R[39]),
		.new_L135_40(new4_L135_R[40]),
		.new_L135_41(new4_L135_R[41]),
		.new_L135_42(new4_L135_R[42]),
		.new_L135_43(new4_L135_R[43]),
		.new_L135_44(new4_L135_R[44]),
		.new_L135_45(new4_L135_R[45]),
		.new_L135_46(new4_L135_R[46]),
		.new_L135_47(new4_L135_R[47]),
		.new_L135_48(new4_L135_R[48]),
		.new_L135_49(new4_L135_R[49]),
		.new_L135_50(new4_L135_R[50]),
		.new_L135_51(new4_L135_R[51]),
		.new_L135_52(new4_L135_R[52]),
		.new_L135_53(new4_L135_R[53]),
		.new_L135_54(new4_L135_R[54]),
		.new_L135_55(new4_L135_R[55]),
		.new_L135_56(new4_L135_R[56]),
		.new_L135_57(new4_L135_R[57]),
		.new_L135_58(new4_L135_R[58]),
		.new_L135_59(new4_L135_R[59]),
		.new_L135_60(new4_L135_R[60]),
		.new_L135_61(new4_L135_R[61]),
		.new_L135_62(new4_L135_R[62]),
		.new_L135_63(new4_L135_R[63]),		
		.en_agg3(en_agg3_R)
		);
	
	agg3#(cost_width) agg3_Right(
		.clk(clk),
		.rst0(rst0_R),
		.rst(rst),
		.clken(clken0),

        .P1(P1),
        .P2(P2),

		.en_first(en_first_R),
		.en_agg3(en_agg3_R),
		.L0_0(new4_L0_R[0]),
		.L0_1(new4_L0_R[1]),
		.L0_2(new4_L0_R[2]),
		.L0_3(new4_L0_R[3]),
		.L0_4(new4_L0_R[4]),
		.L0_5(new4_L0_R[5]),
		.L0_6(new4_L0_R[6]),
		.L0_7(new4_L0_R[7]),
		.L0_8(new4_L0_R[8]),
		.L0_9(new4_L0_R[9]),
		.L0_10(new4_L0_R[10]),
		.L0_11(new4_L0_R[11]),
		.L0_12(new4_L0_R[12]),
		.L0_13(new4_L0_R[13]),
		.L0_14(new4_L0_R[14]),
		.L0_15(new4_L0_R[15]),
		.L0_16(new4_L0_R[16]),
		.L0_17(new4_L0_R[17]),
		.L0_18(new4_L0_R[18]),
		.L0_19(new4_L0_R[19]),
		.L0_20(new4_L0_R[20]),
		.L0_21(new4_L0_R[21]),
		.L0_22(new4_L0_R[22]),
		.L0_23(new4_L0_R[23]),
		.L0_24(new4_L0_R[24]),
		.L0_25(new4_L0_R[25]),
		.L0_26(new4_L0_R[26]),
		.L0_27(new4_L0_R[27]),
		.L0_28(new4_L0_R[28]),
		.L0_29(new4_L0_R[29]),
		.L0_30(new4_L0_R[30]),
		.L0_31(new4_L0_R[31]),
		.L0_32(new4_L0_R[32]),
		.L0_33(new4_L0_R[33]),
		.L0_34(new4_L0_R[34]),
		.L0_35(new4_L0_R[35]),
		.L0_36(new4_L0_R[36]),
		.L0_37(new4_L0_R[37]),
		.L0_38(new4_L0_R[38]),
		.L0_39(new4_L0_R[39]),
		.L0_40(new4_L0_R[40]),
		.L0_41(new4_L0_R[41]),
		.L0_42(new4_L0_R[42]),
		.L0_43(new4_L0_R[43]),
		.L0_44(new4_L0_R[44]),
		.L0_45(new4_L0_R[45]),
		.L0_46(new4_L0_R[46]),
		.L0_47(new4_L0_R[47]),
		.L0_48(new4_L0_R[48]),
		.L0_49(new4_L0_R[49]),
		.L0_50(new4_L0_R[50]),
		.L0_51(new4_L0_R[51]),
		.L0_52(new4_L0_R[52]),
		.L0_53(new4_L0_R[53]),
		.L0_54(new4_L0_R[54]),
		.L0_55(new4_L0_R[55]),
		.L0_56(new4_L0_R[56]),
		.L0_57(new4_L0_R[57]),
		.L0_58(new4_L0_R[58]),
		.L0_59(new4_L0_R[59]),
		.L0_60(new4_L0_R[60]),
		.L0_61(new4_L0_R[61]),
		.L0_62(new4_L0_R[62]),
		.L0_63(new4_L0_R[63]),
		
		.L135_0(new4_L135_R[0]),
		.L135_1(new4_L135_R[1]),
		.L135_2(new4_L135_R[2]),
		.L135_3(new4_L135_R[3]),
		.L135_4(new4_L135_R[4]),
		.L135_5(new4_L135_R[5]),
		.L135_6(new4_L135_R[6]),
		.L135_7(new4_L135_R[7]),
		.L135_8(new4_L135_R[8]),
		.L135_9(new4_L135_R[9]),
		.L135_10(new4_L135_R[10]),
		.L135_11(new4_L135_R[11]),
		.L135_12(new4_L135_R[12]),
		.L135_13(new4_L135_R[13]),
		.L135_14(new4_L135_R[14]),
		.L135_15(new4_L135_R[15]),
		.L135_16(new4_L135_R[16]),
		.L135_17(new4_L135_R[17]),
		.L135_18(new4_L135_R[18]),
		.L135_19(new4_L135_R[19]),
		.L135_20(new4_L135_R[20]),
		.L135_21(new4_L135_R[21]),
		.L135_22(new4_L135_R[22]),
		.L135_23(new4_L135_R[23]),
		.L135_24(new4_L135_R[24]),
		.L135_25(new4_L135_R[25]),
		.L135_26(new4_L135_R[26]),
		.L135_27(new4_L135_R[27]),
		.L135_28(new4_L135_R[28]),
		.L135_29(new4_L135_R[29]),
		.L135_30(new4_L135_R[30]),
		.L135_31(new4_L135_R[31]),
		.L135_32(new4_L135_R[32]),
		.L135_33(new4_L135_R[33]),
		.L135_34(new4_L135_R[34]),
		.L135_35(new4_L135_R[35]),
		.L135_36(new4_L135_R[36]),
		.L135_37(new4_L135_R[37]),
		.L135_38(new4_L135_R[38]),
		.L135_39(new4_L135_R[39]),
		.L135_40(new4_L135_R[40]),
		.L135_41(new4_L135_R[41]),
		.L135_42(new4_L135_R[42]),
		.L135_43(new4_L135_R[43]),
		.L135_44(new4_L135_R[44]),
		.L135_45(new4_L135_R[45]),
		.L135_46(new4_L135_R[46]),
		.L135_47(new4_L135_R[47]),
		.L135_48(new4_L135_R[48]),
		.L135_49(new4_L135_R[49]),
		.L135_50(new4_L135_R[50]),
		.L135_51(new4_L135_R[51]),
		.L135_52(new4_L135_R[52]),
		.L135_53(new4_L135_R[53]),
		.L135_54(new4_L135_R[54]),
		.L135_55(new4_L135_R[55]),
		.L135_56(new4_L135_R[56]),
		.L135_57(new4_L135_R[57]),
		.L135_58(new4_L135_R[58]),
		.L135_59(new4_L135_R[59]),
		.L135_60(new4_L135_R[60]),
		.L135_61(new4_L135_R[61]),
		.L135_62(new4_L135_R[62]),
		.L135_63(new4_L135_R[63]),
		
		.min_135(min_135_R),
	
		.agg135_0(L_135_R[0][2]),
		.agg135_1(L_135_R[1][2]),
		.agg135_2(L_135_R[2][2]),
		.agg135_3(L_135_R[3][2]),
		.agg135_4(L_135_R[4][2]),
		.agg135_5(L_135_R[5][2]),
		.agg135_6(L_135_R[6][2]),
		.agg135_7(L_135_R[7][2]),
		.agg135_8(L_135_R[8][2]),
		.agg135_9(L_135_R[9][2]),
		.agg135_10(L_135_R[10][2]),
		.agg135_11(L_135_R[11][2]),
		.agg135_12(L_135_R[12][2]),
		.agg135_13(L_135_R[13][2]),
		.agg135_14(L_135_R[14][2]),
		.agg135_15(L_135_R[15][2]),
		.agg135_16(L_135_R[16][2]),
		.agg135_17(L_135_R[17][2]),
		.agg135_18(L_135_R[18][2]),
		.agg135_19(L_135_R[19][2]),
		.agg135_20(L_135_R[20][2]),
		.agg135_21(L_135_R[21][2]),
		.agg135_22(L_135_R[22][2]),
		.agg135_23(L_135_R[23][2]),
		.agg135_24(L_135_R[24][2]),
		.agg135_25(L_135_R[25][2]),
		.agg135_26(L_135_R[26][2]),
		.agg135_27(L_135_R[27][2]),
		.agg135_28(L_135_R[28][2]),
		.agg135_29(L_135_R[29][2]),
		.agg135_30(L_135_R[30][2]),
		.agg135_31(L_135_R[31][2]),
		.agg135_32(L_135_R[32][2]),
		.agg135_33(L_135_R[33][2]),
		.agg135_34(L_135_R[34][2]),
		.agg135_35(L_135_R[35][2]),
		.agg135_36(L_135_R[36][2]),
		.agg135_37(L_135_R[37][2]),
		.agg135_38(L_135_R[38][2]),
		.agg135_39(L_135_R[39][2]),
		.agg135_40(L_135_R[40][2]),
		.agg135_41(L_135_R[41][2]),
		.agg135_42(L_135_R[42][2]),
		.agg135_43(L_135_R[43][2]),
		.agg135_44(L_135_R[44][2]),
		.agg135_45(L_135_R[45][2]),
		.agg135_46(L_135_R[46][2]),
		.agg135_47(L_135_R[47][2]),
		.agg135_48(L_135_R[48][2]),
		.agg135_49(L_135_R[49][2]),
		.agg135_50(L_135_R[50][2]),
		.agg135_51(L_135_R[51][2]),
		.agg135_52(L_135_R[52][2]),
		.agg135_53(L_135_R[53][2]),
		.agg135_54(L_135_R[54][2]),
		.agg135_55(L_135_R[55][2]),
		.agg135_56(L_135_R[56][2]),
		.agg135_57(L_135_R[57][2]),
		.agg135_58(L_135_R[58][2]),
		.agg135_59(L_135_R[59][2]),
		.agg135_60(L_135_R[60][2]),
		.agg135_61(L_135_R[61][2]),	
		.agg135_62(L_135_R[62][2]),
		.agg135_63(L_135_R[63][2]),
		
		.new_L0_0(new3_L0_R[0]),
		.new_L0_1(new3_L0_R[1]),
		.new_L0_2(new3_L0_R[2]),
		.new_L0_3(new3_L0_R[3]),
		.new_L0_4(new3_L0_R[4]),
		.new_L0_5(new3_L0_R[5]),
		.new_L0_6(new3_L0_R[6]),
		.new_L0_7(new3_L0_R[7]),
		.new_L0_8(new3_L0_R[8]),
		.new_L0_9(new3_L0_R[9]),
		.new_L0_10(new3_L0_R[10]),
		.new_L0_11(new3_L0_R[11]),
		.new_L0_12(new3_L0_R[12]),
		.new_L0_13(new3_L0_R[13]),
		.new_L0_14(new3_L0_R[14]),
		.new_L0_15(new3_L0_R[15]),
		.new_L0_16(new3_L0_R[16]),
		.new_L0_17(new3_L0_R[17]),
		.new_L0_18(new3_L0_R[18]),
		.new_L0_19(new3_L0_R[19]),
		.new_L0_20(new3_L0_R[20]),
		.new_L0_21(new3_L0_R[21]),
		.new_L0_22(new3_L0_R[22]),
		.new_L0_23(new3_L0_R[23]),
		.new_L0_24(new3_L0_R[24]),
		.new_L0_25(new3_L0_R[25]),
		.new_L0_26(new3_L0_R[26]),
		.new_L0_27(new3_L0_R[27]),
		.new_L0_28(new3_L0_R[28]),
		.new_L0_29(new3_L0_R[29]),
		.new_L0_30(new3_L0_R[30]),
		.new_L0_31(new3_L0_R[31]),
		.new_L0_32(new3_L0_R[32]),
		.new_L0_33(new3_L0_R[33]),
		.new_L0_34(new3_L0_R[34]),
		.new_L0_35(new3_L0_R[35]),
		.new_L0_36(new3_L0_R[36]),
		.new_L0_37(new3_L0_R[37]),
		.new_L0_38(new3_L0_R[38]),
		.new_L0_39(new3_L0_R[39]),
		.new_L0_40(new3_L0_R[40]),
		.new_L0_41(new3_L0_R[41]),
		.new_L0_42(new3_L0_R[42]),
		.new_L0_43(new3_L0_R[43]),
		.new_L0_44(new3_L0_R[44]),
		.new_L0_45(new3_L0_R[45]),
		.new_L0_46(new3_L0_R[46]),
		.new_L0_47(new3_L0_R[47]),
		.new_L0_48(new3_L0_R[48]),
		.new_L0_49(new3_L0_R[49]),
		.new_L0_50(new3_L0_R[50]),
		.new_L0_51(new3_L0_R[51]),
		.new_L0_52(new3_L0_R[52]),
		.new_L0_53(new3_L0_R[53]),
		.new_L0_54(new3_L0_R[54]),
		.new_L0_55(new3_L0_R[55]),
		.new_L0_56(new3_L0_R[56]),
		.new_L0_57(new3_L0_R[57]),
		.new_L0_58(new3_L0_R[58]),
		.new_L0_59(new3_L0_R[59]),
		.new_L0_60(new3_L0_R[60]),
		.new_L0_61(new3_L0_R[61]),
		.new_L0_62(new3_L0_R[62]),
		.new_L0_63(new3_L0_R[63]),
			
		.new_L135_0(new3_L135_R[0]),
		.new_L135_1(new3_L135_R[1]),
		.new_L135_2(new3_L135_R[2]),
		.new_L135_3(new3_L135_R[3]),
		.new_L135_4(new3_L135_R[4]),
		.new_L135_5(new3_L135_R[5]),
		.new_L135_6(new3_L135_R[6]),
		.new_L135_7(new3_L135_R[7]),
		.new_L135_8(new3_L135_R[8]),
		.new_L135_9(new3_L135_R[9]),
		.new_L135_10(new3_L135_R[10]),
		.new_L135_11(new3_L135_R[11]),
		.new_L135_12(new3_L135_R[12]),
		.new_L135_13(new3_L135_R[13]),
		.new_L135_14(new3_L135_R[14]),
		.new_L135_15(new3_L135_R[15]),
		.new_L135_16(new3_L135_R[16]),
		.new_L135_17(new3_L135_R[17]),
		.new_L135_18(new3_L135_R[18]),
		.new_L135_19(new3_L135_R[19]),
		.new_L135_20(new3_L135_R[20]),
		.new_L135_21(new3_L135_R[21]),
		.new_L135_22(new3_L135_R[22]),
		.new_L135_23(new3_L135_R[23]),
		.new_L135_24(new3_L135_R[24]),
		.new_L135_25(new3_L135_R[25]),
		.new_L135_26(new3_L135_R[26]),
		.new_L135_27(new3_L135_R[27]),
		.new_L135_28(new3_L135_R[28]),
		.new_L135_29(new3_L135_R[29]),
		.new_L135_30(new3_L135_R[30]),
		.new_L135_31(new3_L135_R[31]),
		.new_L135_32(new3_L135_R[32]),
		.new_L135_33(new3_L135_R[33]),
		.new_L135_34(new3_L135_R[34]),
		.new_L135_35(new3_L135_R[35]),
		.new_L135_36(new3_L135_R[36]),
		.new_L135_37(new3_L135_R[37]),
		.new_L135_38(new3_L135_R[38]),
		.new_L135_39(new3_L135_R[39]),
		.new_L135_40(new3_L135_R[40]),
		.new_L135_41(new3_L135_R[41]),
		.new_L135_42(new3_L135_R[42]),
		.new_L135_43(new3_L135_R[43]),
		.new_L135_44(new3_L135_R[44]),
		.new_L135_45(new3_L135_R[45]),
		.new_L135_46(new3_L135_R[46]),
		.new_L135_47(new3_L135_R[47]),
		.new_L135_48(new3_L135_R[48]),
		.new_L135_49(new3_L135_R[49]),
		.new_L135_50(new3_L135_R[50]),
		.new_L135_51(new3_L135_R[51]),
		.new_L135_52(new3_L135_R[52]),
		.new_L135_53(new3_L135_R[53]),
		.new_L135_54(new3_L135_R[54]),
		.new_L135_55(new3_L135_R[55]),
		.new_L135_56(new3_L135_R[56]),
		.new_L135_57(new3_L135_R[57]),
		.new_L135_58(new3_L135_R[58]),
		.new_L135_59(new3_L135_R[59]),
		.new_L135_60(new3_L135_R[60]),
		.new_L135_61(new3_L135_R[61]),
		.new_L135_62(new3_L135_R[62]),
		.new_L135_63(new3_L135_R[63]),
	
		.en_disp(en_disp_R),
	
		.cost_valid(cost_valid)
		);
		//disparity for the right direction
	
	disparity#(cost_width)  disparity_Right(
	
			.rst(rst),
	
			.clk(clk),
	
			.clken(clken0),
	
			.en_disp(en_agg3_R),
	
			//0?
			.aggregateCost0_0(L_0_R[0][2]),
			.aggregateCost0_1(L_0_R[1][2]),
			.aggregateCost0_2(L_0_R[2][2]), 
			.aggregateCost0_3(L_0_R[3][2]),
			.aggregateCost0_4(L_0_R[4][2]),
			.aggregateCost0_5(L_0_R[5][2]), 
			.aggregateCost0_6(L_0_R[6][2]),
			.aggregateCost0_7(L_0_R[7][2]),
			.aggregateCost0_8(L_0_R[8][2]), 
			.aggregateCost0_9(L_0_R[9][2]),
			.aggregateCost0_10(L_0_R[10][2]),
			.aggregateCost0_11(L_0_R[11][2]), 
			.aggregateCost0_12(L_0_R[12][2]),
			.aggregateCost0_13(L_0_R[13][2]),
			.aggregateCost0_14(L_0_R[14][2]), 
			.aggregateCost0_15(L_0_R[15][2]),
			.aggregateCost0_16(L_0_R[16][2]),
			.aggregateCost0_17(L_0_R[17][2]), 
			.aggregateCost0_18(L_0_R[18][2]),
			.aggregateCost0_19(L_0_R[19][2]),
			.aggregateCost0_20(L_0_R[20][2]), 
			.aggregateCost0_21(L_0_R[21][2]),
			.aggregateCost0_22(L_0_R[22][2]),
			.aggregateCost0_23(L_0_R[23][2]), 
			.aggregateCost0_24(L_0_R[24][2]), 
			.aggregateCost0_25(L_0_R[25][2]),
			.aggregateCost0_26(L_0_R[26][2]),
			.aggregateCost0_27(L_0_R[27][2]), 
			.aggregateCost0_28(L_0_R[28][2]), 
			.aggregateCost0_29(L_0_R[29][2]),
			.aggregateCost0_30(L_0_R[30][2]),
			.aggregateCost0_31(L_0_R[31][2]), 
			.aggregateCost0_32(L_0_R[32][2]), 
			.aggregateCost0_33(L_0_R[33][2]),
			.aggregateCost0_34(L_0_R[34][2]),
			.aggregateCost0_35(L_0_R[35][2]), 
			.aggregateCost0_36(L_0_R[36][2]),
			.aggregateCost0_37(L_0_R[37][2]),
			.aggregateCost0_38(L_0_R[38][2]), 
			.aggregateCost0_39(L_0_R[39][2]),
			.aggregateCost0_40(L_0_R[40][2]),
			.aggregateCost0_41(L_0_R[41][2]), 
			.aggregateCost0_42(L_0_R[42][2]),
			.aggregateCost0_43(L_0_R[43][2]),
			.aggregateCost0_44(L_0_R[44][2]), 
			.aggregateCost0_45(L_0_R[45][2]),
			.aggregateCost0_46(L_0_R[46][2]),
			.aggregateCost0_47(L_0_R[47][2]), 
			.aggregateCost0_48(L_0_R[48][2]),
			.aggregateCost0_49(L_0_R[49][2]),
			.aggregateCost0_50(L_0_R[50][2]), 
			.aggregateCost0_51(L_0_R[51][2]),
			.aggregateCost0_52(L_0_R[52][2]),
			.aggregateCost0_53(L_0_R[53][2]), 
			.aggregateCost0_54(L_0_R[54][2]), 
			.aggregateCost0_55(L_0_R[55][2]),
			.aggregateCost0_56(L_0_R[56][2]),
			.aggregateCost0_57(L_0_R[57][2]), 
			.aggregateCost0_58(L_0_R[58][2]), 
			.aggregateCost0_59(L_0_R[59][2]),
			.aggregateCost0_60(L_0_R[60][2]),
			.aggregateCost0_61(L_0_R[61][2]),
			.aggregateCost0_62(L_0_R[62][2]),
			.aggregateCost0_63(L_0_R[63][2]),		
	
			//135?
			.aggregateCost3_0(L_135_R[0][2]),
			.aggregateCost3_1(L_135_R[1][2]),
			.aggregateCost3_2(L_135_R[2][2]), 
			.aggregateCost3_3(L_135_R[3][2]),
			.aggregateCost3_4(L_135_R[4][2]),
			.aggregateCost3_5(L_135_R[5][2]), 
			.aggregateCost3_6(L_135_R[6][2]),
			.aggregateCost3_7(L_135_R[7][2]),
			.aggregateCost3_8(L_135_R[8][2]), 
			.aggregateCost3_9(L_135_R[9][2]),
			.aggregateCost3_10(L_135_R[10][2]),
			.aggregateCost3_11(L_135_R[11][2]), 
			.aggregateCost3_12(L_135_R[12][2]),
			.aggregateCost3_13(L_135_R[13][2]),
			.aggregateCost3_14(L_135_R[14][2]), 
			.aggregateCost3_15(L_135_R[15][2]),
			.aggregateCost3_16(L_135_R[16][2]),
			.aggregateCost3_17(L_135_R[17][2]), 
			.aggregateCost3_18(L_135_R[18][2]),
			.aggregateCost3_19(L_135_R[19][2]),
			.aggregateCost3_20(L_135_R[20][2]), 
			.aggregateCost3_21(L_135_R[21][2]),
			.aggregateCost3_22(L_135_R[22][2]),
			.aggregateCost3_23(L_135_R[23][2]), 
			.aggregateCost3_24(L_135_R[24][2]), 
			.aggregateCost3_25(L_135_R[25][2]),
			.aggregateCost3_26(L_135_R[26][2]),
			.aggregateCost3_27(L_135_R[27][2]), 
			.aggregateCost3_28(L_135_R[28][2]), 
			.aggregateCost3_29(L_135_R[29][2]),
			.aggregateCost3_30(L_135_R[30][2]),
			.aggregateCost3_31(L_135_R[31][2]), 
			.aggregateCost3_32(L_135_R[32][2]), 
			.aggregateCost3_33(L_135_R[33][2]),
			.aggregateCost3_34(L_135_R[34][2]),
			.aggregateCost3_35(L_135_R[35][2]), 
			.aggregateCost3_36(L_135_R[36][2]),
			.aggregateCost3_37(L_135_R[37][2]),
			.aggregateCost3_38(L_135_R[38][2]), 
			.aggregateCost3_39(L_135_R[39][2]),
			.aggregateCost3_40(L_135_R[40][2]),
			.aggregateCost3_41(L_135_R[41][2]), 
			.aggregateCost3_42(L_135_R[42][2]),
			.aggregateCost3_43(L_135_R[43][2]),
			.aggregateCost3_44(L_135_R[44][2]), 
			.aggregateCost3_45(L_135_R[45][2]),
			.aggregateCost3_46(L_135_R[46][2]),
			.aggregateCost3_47(L_135_R[47][2]), 
			.aggregateCost3_48(L_135_R[48][2]),
			.aggregateCost3_49(L_135_R[49][2]),
			.aggregateCost3_50(L_135_R[50][2]), 
			.aggregateCost3_51(L_135_R[51][2]),
			.aggregateCost3_52(L_135_R[52][2]),
			.aggregateCost3_53(L_135_R[53][2]), 
			.aggregateCost3_54(L_135_R[54][2]), 
			.aggregateCost3_55(L_135_R[55][2]),
			.aggregateCost3_56(L_135_R[56][2]),
			.aggregateCost3_57(L_135_R[57][2]), 
			.aggregateCost3_58(L_135_R[58][2]), 
			.aggregateCost3_59(L_135_R[59][2]),
			.aggregateCost3_60(L_135_R[60][2]),
			.aggregateCost3_61(L_135_R[61][2]),
			.aggregateCost3_62(L_135_R[62][2]),
			.aggregateCost3_63(L_135_R[63][2]),
	
			.disp_final(disp_R),
	
			.valid_final(valid_final_R),
			
			.cost_valid(cost_valid)
	
			);
	
		
	
	
	
	
	
	//left
	wire  [cost_width-1:0] min_0_L;
	
	
	reg en_first_L;
	reg en_first_L_agg2;
	wire en_agg3_L;
	
	
	wire  [cost_width-3:0] min_135_L;
	
	//agg3
	wire en_disp_L;
	wire valid_1_L;	
	wire valid_2_L;
	reg change_L;
	wire valid_3_L;
	//middle
	wire  [cost_width-1:0]L_0_L[63:0][2:0];
	wire  [cost_width-3:0]L_135_L[63:0][2:0];
	
	wire [cost_width-1:0] new3_L0_L[63:0];
	wire [cost_width-3:0] new3_L135_L[63:0];
	wire [cost_width-1:0] L_3_0_L[63:0];
	wire [cost_width-3:0] L_3_135_L[63:0];
	
	assign L_0_L[0][0]=L_3_0_L[0];
	assign L_0_L[1][0]=L_3_0_L[1];
	assign L_0_L[2][0]=L_3_0_L[2];
	assign L_0_L[3][0]=L_3_0_L[3];
	assign L_0_L[4][0]=L_3_0_L[4];
	assign L_0_L[5][0]=L_3_0_L[5];
	assign L_0_L[6][0]=L_3_0_L[6];
	assign L_0_L[7][0]=L_3_0_L[7];
	assign L_0_L[8][0]=L_3_0_L[8];
	assign L_0_L[9][0]=L_3_0_L[9];
	assign L_0_L[10][0]=L_3_0_L[10];
	assign L_0_L[11][0]=L_3_0_L[11];
	assign L_0_L[12][0]=L_3_0_L[12];
	assign L_0_L[13][0]=L_3_0_L[13];
	assign L_0_L[14][0]=L_3_0_L[14];
	assign L_0_L[15][0]=L_3_0_L[15];
	assign L_0_L[16][0]=L_3_0_L[16];
	assign L_0_L[17][0]=L_3_0_L[17];
	assign L_0_L[18][0]=L_3_0_L[18];
	assign L_0_L[19][0]=L_3_0_L[19];
	assign L_0_L[20][0]=L_3_0_L[20];
	assign L_0_L[21][0]=L_3_0_L[21];
	assign L_0_L[22][0]=L_3_0_L[22];
	assign L_0_L[23][0]=L_3_0_L[23];
	assign L_0_L[24][0]=L_3_0_L[24];
	assign L_0_L[25][0]=L_3_0_L[25];
	assign L_0_L[26][0]=L_3_0_L[26];
	assign L_0_L[27][0]=L_3_0_L[27];
	assign L_0_L[28][0]=L_3_0_L[28];
	assign L_0_L[29][0]=L_3_0_L[29];
	assign L_0_L[30][0]=L_3_0_L[30];
	assign L_0_L[31][0]=L_3_0_L[31];
	assign L_0_L[32][0]=L_3_0_L[32];
	assign L_0_L[33][0]=L_3_0_L[33];
	assign L_0_L[34][0]=L_3_0_L[34];
	assign L_0_L[35][0]=L_3_0_L[35];
	assign L_0_L[36][0]=L_3_0_L[36];
	assign L_0_L[37][0]=L_3_0_L[37];
	assign L_0_L[38][0]=L_3_0_L[38];
	assign L_0_L[39][0]=L_3_0_L[39];
	assign L_0_L[40][0]=L_3_0_L[40];
	assign L_0_L[41][0]=L_3_0_L[41];
	assign L_0_L[42][0]=L_3_0_L[42];
	assign L_0_L[43][0]=L_3_0_L[43];
	assign L_0_L[44][0]=L_3_0_L[44];
	assign L_0_L[45][0]=L_3_0_L[45];
	assign L_0_L[46][0]=L_3_0_L[46];
	assign L_0_L[47][0]=L_3_0_L[47];
	assign L_0_L[48][0]=L_3_0_L[48];
	assign L_0_L[49][0]=L_3_0_L[49];
	assign L_0_L[50][0]=L_3_0_L[50];
	assign L_0_L[51][0]=L_3_0_L[51];
	assign L_0_L[52][0]=L_3_0_L[52];
	assign L_0_L[53][0]=L_3_0_L[53];
	assign L_0_L[54][0]=L_3_0_L[54];
	assign L_0_L[55][0]=L_3_0_L[55];
	assign L_0_L[56][0]=L_3_0_L[56];
	assign L_0_L[57][0]=L_3_0_L[57];
	assign L_0_L[58][0]=L_3_0_L[58];
	assign L_0_L[59][0]=L_3_0_L[59];
	assign L_0_L[60][0]=L_3_0_L[60];
	assign L_0_L[61][0]=L_3_0_L[61];
	assign L_0_L[62][0]=L_3_0_L[62];
	assign L_0_L[63][0]=L_3_0_L[63];
	
	assign L_135_L[0][0]=L_3_135_L[0];
	assign L_135_L[1][0]=L_3_135_L[1];
	assign L_135_L[2][0]=L_3_135_L[2];
	assign L_135_L[3][0]=L_3_135_L[3];
	assign L_135_L[4][0]=L_3_135_L[4];
	assign L_135_L[5][0]=L_3_135_L[5];
	assign L_135_L[6][0]=L_3_135_L[6];
	assign L_135_L[7][0]=L_3_135_L[7];
	assign L_135_L[8][0]=L_3_135_L[8];
	assign L_135_L[9][0]=L_3_135_L[9];
	assign L_135_L[10][0]=L_3_135_L[10];
	assign L_135_L[11][0]=L_3_135_L[11];
	assign L_135_L[12][0]=L_3_135_L[12];
	assign L_135_L[13][0]=L_3_135_L[13];
	assign L_135_L[14][0]=L_3_135_L[14];
	assign L_135_L[15][0]=L_3_135_L[15];
	assign L_135_L[16][0]=L_3_135_L[16];
	assign L_135_L[17][0]=L_3_135_L[17];
	assign L_135_L[18][0]=L_3_135_L[18];
	assign L_135_L[19][0]=L_3_135_L[19];
	assign L_135_L[20][0]=L_3_135_L[20];
	assign L_135_L[21][0]=L_3_135_L[21];
	assign L_135_L[22][0]=L_3_135_L[22];
	assign L_135_L[23][0]=L_3_135_L[23];
	assign L_135_L[24][0]=L_3_135_L[24];
	assign L_135_L[25][0]=L_3_135_L[25];
	assign L_135_L[26][0]=L_3_135_L[26];
	assign L_135_L[27][0]=L_3_135_L[27];
	assign L_135_L[28][0]=L_3_135_L[28];
	assign L_135_L[29][0]=L_3_135_L[29];
	assign L_135_L[30][0]=L_3_135_L[30];
	assign L_135_L[31][0]=L_3_135_L[31];
	assign L_135_L[32][0]=L_3_135_L[32];
	assign L_135_L[33][0]=L_3_135_L[33];
	assign L_135_L[34][0]=L_3_135_L[34];
	assign L_135_L[35][0]=L_3_135_L[35];
	assign L_135_L[36][0]=L_3_135_L[36];
	assign L_135_L[37][0]=L_3_135_L[37];
	assign L_135_L[38][0]=L_3_135_L[38];
	assign L_135_L[39][0]=L_3_135_L[39];
	assign L_135_L[40][0]=L_3_135_L[40];
	assign L_135_L[41][0]=L_3_135_L[41];
	assign L_135_L[42][0]=L_3_135_L[42];
	assign L_135_L[43][0]=L_3_135_L[43];
	assign L_135_L[44][0]=L_3_135_L[44];
	assign L_135_L[45][0]=L_3_135_L[45];
	assign L_135_L[46][0]=L_3_135_L[46];
	assign L_135_L[47][0]=L_3_135_L[47];
	assign L_135_L[48][0]=L_3_135_L[48];
	assign L_135_L[49][0]=L_3_135_L[49];
	assign L_135_L[50][0]=L_3_135_L[50];
	assign L_135_L[51][0]=L_3_135_L[51];
	assign L_135_L[52][0]=L_3_135_L[52];
	assign L_135_L[53][0]=L_3_135_L[53];
	assign L_135_L[54][0]=L_3_135_L[54];
	assign L_135_L[55][0]=L_3_135_L[55];
	assign L_135_L[56][0]=L_3_135_L[56];
	assign L_135_L[57][0]=L_3_135_L[57];
	assign L_135_L[58][0]=L_3_135_L[58];
	assign L_135_L[59][0]=L_3_135_L[59];
	assign L_135_L[60][0]=L_3_135_L[60];
	assign L_135_L[61][0]=L_3_135_L[61];
	assign L_135_L[62][0]=L_3_135_L[62];
	assign L_135_L[63][0]=L_3_135_L[63];
	
	reg en_agg4_L;
	reg rst0_L;	
	
	wire [cost_width-1:0] L0_L[63:0];
	wire [cost_width-3:0] L135_L[63:0];
	
	agg_first#(cost_width) agg_first_Left(
		.clk(clk),
		.rst(rst),
		.clken(clken0),
		.valid(en_L),
		.valid_1(valid_1_L),
		
		.cost0_0(cost_L_in[0]),
		.cost0_1(cost_L_in[1]),
		.cost0_2(cost_L_in[2]),
		.cost0_3(cost_L_in[3]),
		.cost0_4(cost_L_in[4]),
		.cost0_5(cost_L_in[5]),
		.cost0_6(cost_L_in[6]),
		.cost0_7(cost_L_in[7]),
		.cost0_8(cost_L_in[8]),
		.cost0_9(cost_L_in[9]),
		.cost0_10(cost_L_in[10]),
		.cost0_11(cost_L_in[11]),
		.cost0_12(cost_L_in[12]),
		.cost0_13(cost_L_in[13]),
		.cost0_14(cost_L_in[14]),
		.cost0_15(cost_L_in[15]),
		.cost0_16(cost_L_in[16]),
		.cost0_17(cost_L_in[17]),
		.cost0_18(cost_L_in[18]),
		.cost0_19(cost_L_in[19]),
		.cost0_20(cost_L_in[20]),
		.cost0_21(cost_L_in[21]),
		.cost0_22(cost_L_in[22]),
		.cost0_23(cost_L_in[23]),
		.cost0_24(cost_L_in[24]),
		.cost0_25(cost_L_in[25]),
		.cost0_26(cost_L_in[26]),
		.cost0_27(cost_L_in[27]),
		.cost0_28(cost_L_in[28]),
		.cost0_29(cost_L_in[29]),
		.cost0_30(cost_L_in[30]),
		.cost0_31(cost_L_in[31]),
		.cost0_32(cost_L_in[32]),
		.cost0_33(cost_L_in[33]),
		.cost0_34(cost_L_in[34]),
		.cost0_35(cost_L_in[35]),
		.cost0_36(cost_L_in[36]),
		.cost0_37(cost_L_in[37]),
		.cost0_38(cost_L_in[38]),
		.cost0_39(cost_L_in[39]),
		.cost0_40(cost_L_in[40]),
		.cost0_41(cost_L_in[41]),
		.cost0_42(cost_L_in[42]),
		.cost0_43(cost_L_in[43]),
		.cost0_44(cost_L_in[44]),
		.cost0_45(cost_L_in[45]),
		.cost0_46(cost_L_in[46]),
		.cost0_47(cost_L_in[47]),
		.cost0_48(cost_L_in[48]),
		.cost0_49(cost_L_in[49]),
		.cost0_50(cost_L_in[50]),
		.cost0_51(cost_L_in[51]),
		.cost0_52(cost_L_in[52]),
		.cost0_53(cost_L_in[53]),
		.cost0_54(cost_L_in[54]),
		.cost0_55(cost_L_in[55]),
		.cost0_56(cost_L_in[56]),
		.cost0_57(cost_L_in[57]),
		.cost0_58(cost_L_in[58]),
		.cost0_59(cost_L_in[59]),
		.cost0_60(cost_L_in[60]),
		.cost0_61(cost_L_in[61]),
		.cost0_62(cost_L_in[62]),
		.cost0_63(cost_L_in[63]),
		
		.cost135_0(cost_L_in[0][cost_width-1:2]),
		.cost135_1(cost_L_in[1][cost_width-1:2]),
		.cost135_2(cost_L_in[2][cost_width-1:2]),
		.cost135_3(cost_L_in[3][cost_width-1:2]),
		.cost135_4(cost_L_in[4][cost_width-1:2]),
		.cost135_5(cost_L_in[5][cost_width-1:2]),
		.cost135_6(cost_L_in[6][cost_width-1:2]),
		.cost135_7(cost_L_in[7][cost_width-1:2]),
		.cost135_8(cost_L_in[8][cost_width-1:2]),
		.cost135_9(cost_L_in[9][cost_width-1:2]),
		.cost135_10(cost_L_in[10][cost_width-1:2]),
		.cost135_11(cost_L_in[11][cost_width-1:2]),
		.cost135_12(cost_L_in[12][cost_width-1:2]),
		.cost135_13(cost_L_in[13][cost_width-1:2]),
		.cost135_14(cost_L_in[14][cost_width-1:2]),
		.cost135_15(cost_L_in[15][cost_width-1:2]),
		.cost135_16(cost_L_in[16][cost_width-1:2]),
		.cost135_17(cost_L_in[17][cost_width-1:2]),
		.cost135_18(cost_L_in[18][cost_width-1:2]),
		.cost135_19(cost_L_in[19][cost_width-1:2]),
		.cost135_20(cost_L_in[20][cost_width-1:2]),
		.cost135_21(cost_L_in[21][cost_width-1:2]),
		.cost135_22(cost_L_in[22][cost_width-1:2]),
		.cost135_23(cost_L_in[23][cost_width-1:2]),
		.cost135_24(cost_L_in[24][cost_width-1:2]),
		.cost135_25(cost_L_in[25][cost_width-1:2]),
		.cost135_26(cost_L_in[26][cost_width-1:2]),
		.cost135_27(cost_L_in[27][cost_width-1:2]),
		.cost135_28(cost_L_in[28][cost_width-1:2]),
		.cost135_29(cost_L_in[29][cost_width-1:2]),
		.cost135_30(cost_L_in[30][cost_width-1:2]),
		.cost135_31(cost_L_in[31][cost_width-1:2]),
		.cost135_32(cost_L_in[32][cost_width-1:2]),
		.cost135_33(cost_L_in[33][cost_width-1:2]),
		.cost135_34(cost_L_in[34][cost_width-1:2]),
		.cost135_35(cost_L_in[35][cost_width-1:2]),
		.cost135_36(cost_L_in[36][cost_width-1:2]),
		.cost135_37(cost_L_in[37][cost_width-1:2]),
		.cost135_38(cost_L_in[38][cost_width-1:2]),
		.cost135_39(cost_L_in[39][cost_width-1:2]),
		.cost135_40(cost_L_in[40][cost_width-1:2]),
		.cost135_41(cost_L_in[41][cost_width-1:2]),
		.cost135_42(cost_L_in[42][cost_width-1:2]),
		.cost135_43(cost_L_in[43][cost_width-1:2]),
		.cost135_44(cost_L_in[44][cost_width-1:2]),
		.cost135_45(cost_L_in[45][cost_width-1:2]),
		.cost135_46(cost_L_in[46][cost_width-1:2]),
		.cost135_47(cost_L_in[47][cost_width-1:2]),
		.cost135_48(cost_L_in[48][cost_width-1:2]),
		.cost135_49(cost_L_in[49][cost_width-1:2]),
		.cost135_50(cost_L_in[50][cost_width-1:2]),
		.cost135_51(cost_L_in[51][cost_width-1:2]),
		.cost135_52(cost_L_in[52][cost_width-1:2]),
		.cost135_53(cost_L_in[53][cost_width-1:2]),
		.cost135_54(cost_L_in[54][cost_width-1:2]),
		.cost135_55(cost_L_in[55][cost_width-1:2]),
		.cost135_56(cost_L_in[56][cost_width-1:2]),
		.cost135_57(cost_L_in[57][cost_width-1:2]),
		.cost135_58(cost_L_in[58][cost_width-1:2]),
		.cost135_59(cost_L_in[59][cost_width-1:2]),
		.cost135_60(cost_L_in[60][cost_width-1:2]),
		.cost135_61(cost_L_in[61][cost_width-1:2]),
		.cost135_62(cost_L_in[62][cost_width-1:2]),
		.cost135_63(cost_L_in[63][cost_width-1:2]),
		
		.L0_0(L0_L[0]),
		.L0_1(L0_L[1]),
		.L0_2(L0_L[2]),
		.L0_3(L0_L[3]),
		.L0_4(L0_L[4]),
		.L0_5(L0_L[5]),
		.L0_6(L0_L[6]),
		.L0_7(L0_L[7]),
		.L0_8(L0_L[8]),
		.L0_9(L0_L[9]),
		.L0_10(L0_L[10]),
		.L0_11(L0_L[11]),
		.L0_12(L0_L[12]),
		.L0_13(L0_L[13]),
		.L0_14(L0_L[14]),
		.L0_15(L0_L[15]),
		.L0_16(L0_L[16]),
		.L0_17(L0_L[17]),
		.L0_18(L0_L[18]),
		.L0_19(L0_L[19]),
		.L0_20(L0_L[20]),
		.L0_21(L0_L[21]),
		.L0_22(L0_L[22]),
		.L0_23(L0_L[23]),
		.L0_24(L0_L[24]),
		.L0_25(L0_L[25]),
		.L0_26(L0_L[26]),
		.L0_27(L0_L[27]),
		.L0_28(L0_L[28]),
		.L0_29(L0_L[29]),
		.L0_30(L0_L[30]),
		.L0_31(L0_L[31]),
		.L0_32(L0_L[32]),
		.L0_33(L0_L[33]),
		.L0_34(L0_L[34]),
		.L0_35(L0_L[35]),
		.L0_36(L0_L[36]),
		.L0_37(L0_L[37]),
		.L0_38(L0_L[38]),
		.L0_39(L0_L[39]),
		.L0_40(L0_L[40]),
		.L0_41(L0_L[41]),
		.L0_42(L0_L[42]),
		.L0_43(L0_L[43]),
		.L0_44(L0_L[44]),
		.L0_45(L0_L[45]),
		.L0_46(L0_L[46]),
		.L0_47(L0_L[47]),
		.L0_48(L0_L[48]),
		.L0_49(L0_L[49]),
		.L0_50(L0_L[50]),
		.L0_51(L0_L[51]),
		.L0_52(L0_L[52]),
		.L0_53(L0_L[53]),
		.L0_54(L0_L[54]),
		.L0_55(L0_L[55]),
		.L0_56(L0_L[56]),
		.L0_57(L0_L[57]),
		.L0_58(L0_L[58]),
		.L0_59(L0_L[59]),
		.L0_60(L0_L[60]),
		.L0_61(L0_L[61]),
		.L0_62(L0_L[62]),
		.L0_63(L0_L[63]),
		
		.L135_0(L135_L[0]),
		.L135_1(L135_L[1]),
		.L135_2(L135_L[2]),
		.L135_3(L135_L[3]),
		.L135_4(L135_L[4]),
		.L135_5(L135_L[5]),
		.L135_6(L135_L[6]),
		.L135_7(L135_L[7]),
		.L135_8(L135_L[8]),
		.L135_9(L135_L[9]),
		.L135_10(L135_L[10]),
		.L135_11(L135_L[11]),
		.L135_12(L135_L[12]),
		.L135_13(L135_L[13]),
		.L135_14(L135_L[14]),
		.L135_15(L135_L[15]),
		.L135_16(L135_L[16]),
		.L135_17(L135_L[17]),
		.L135_18(L135_L[18]),
		.L135_19(L135_L[19]),
		.L135_20(L135_L[20]),
		.L135_21(L135_L[21]),
		.L135_22(L135_L[22]),
		.L135_23(L135_L[23]),
		.L135_24(L135_L[24]),
		.L135_25(L135_L[25]),
		.L135_26(L135_L[26]),
		.L135_27(L135_L[27]),
		.L135_28(L135_L[28]),
		.L135_29(L135_L[29]),
		.L135_30(L135_L[30]),
		.L135_31(L135_L[31]),
		.L135_32(L135_L[32]),
		.L135_33(L135_L[33]),
		.L135_34(L135_L[34]),
		.L135_35(L135_L[35]),
		.L135_36(L135_L[36]),
		.L135_37(L135_L[37]),
		.L135_38(L135_L[38]),
		.L135_39(L135_L[39]),
		.L135_40(L135_L[40]),
		.L135_41(L135_L[41]),
		.L135_42(L135_L[42]),
		.L135_43(L135_L[43]),
		.L135_44(L135_L[44]),
		.L135_45(L135_L[45]),
		.L135_46(L135_L[46]),
		.L135_47(L135_L[47]),
		.L135_48(L135_L[48]),
		.L135_49(L135_L[49]),
		.L135_50(L135_L[50]),
		.L135_51(L135_L[51]),
		.L135_52(L135_L[52]),
		.L135_53(L135_L[53]),
		.L135_54(L135_L[54]),
		.L135_55(L135_L[55]),
		.L135_56(L135_L[56]),
		.L135_57(L135_L[57]),
		.L135_58(L135_L[58]),
		.L135_59(L135_L[59]),
		.L135_60(L135_L[60]),
		.L135_61(L135_L[61]),
		.L135_62(L135_L[62]),
		.L135_63(L135_L[63])
		
		);
	
	wire [cost_width-1:0] L_2_0_L[63:0];
	wire [cost_width-3:0] L_2_135_L[63:0];
	
	agg_second#(cost_width) agg_second_Left(
		.clk(clk),
		.rst(rst),
		.clken(clken0),
		.valid_1(valid_1_L),
		.valid_2(valid_2_L),
		.cost0_0(L0_L[0]),
		.cost0_1(L0_L[1]),
		.cost0_2(L0_L[2]),
		.cost0_3(L0_L[3]),
		.cost0_4(L0_L[4]),
		.cost0_5(L0_L[5]),
		.cost0_6(L0_L[6]),
		.cost0_7(L0_L[7]),
		.cost0_8(L0_L[8]),
		.cost0_9(L0_L[9]),
		.cost0_10(L0_L[10]),
		.cost0_11(L0_L[11]),
		.cost0_12(L0_L[12]),
		.cost0_13(L0_L[13]),
		.cost0_14(L0_L[14]),
		.cost0_15(L0_L[15]),
		.cost0_16(L0_L[16]),
		.cost0_17(L0_L[17]),
		.cost0_18(L0_L[18]),
		.cost0_19(L0_L[19]),
		.cost0_20(L0_L[20]),
		.cost0_21(L0_L[21]),
		.cost0_22(L0_L[22]),
		.cost0_23(L0_L[23]),
		.cost0_24(L0_L[24]),
		.cost0_25(L0_L[25]),
		.cost0_26(L0_L[26]),
		.cost0_27(L0_L[27]),
		.cost0_28(L0_L[28]),
		.cost0_29(L0_L[29]),
		.cost0_30(L0_L[30]),
		.cost0_31(L0_L[31]),
		.cost0_32(L0_L[32]),
		.cost0_33(L0_L[33]),
		.cost0_34(L0_L[34]),
		.cost0_35(L0_L[35]),
		.cost0_36(L0_L[36]),
		.cost0_37(L0_L[37]),
		.cost0_38(L0_L[38]),
		.cost0_39(L0_L[39]),
		.cost0_40(L0_L[40]),
		.cost0_41(L0_L[41]),
		.cost0_42(L0_L[42]),
		.cost0_43(L0_L[43]),
		.cost0_44(L0_L[44]),
		.cost0_45(L0_L[45]),
		.cost0_46(L0_L[46]),
		.cost0_47(L0_L[47]),
		.cost0_48(L0_L[48]),
		.cost0_49(L0_L[49]),
		.cost0_50(L0_L[50]),
		.cost0_51(L0_L[51]),
		.cost0_52(L0_L[52]),
		.cost0_53(L0_L[53]),
		.cost0_54(L0_L[54]),
		.cost0_55(L0_L[55]),
		.cost0_56(L0_L[56]),
		.cost0_57(L0_L[57]),
		.cost0_58(L0_L[58]),
		.cost0_59(L0_L[59]),
		.cost0_60(L0_L[60]),
		.cost0_61(L0_L[61]),
		.cost0_62(L0_L[62]),
		.cost0_63(L0_L[63]),
	
		.cost135_0(L135_L[0]),
		.cost135_1(L135_L[1]),
		.cost135_2(L135_L[2]),
		.cost135_3(L135_L[3]),
		.cost135_4(L135_L[4]),
		.cost135_5(L135_L[5]),
		.cost135_6(L135_L[6]),
		.cost135_7(L135_L[7]),
		.cost135_8(L135_L[8]),
		.cost135_9(L135_L[9]),
		.cost135_10(L135_L[10]),
		.cost135_11(L135_L[11]),
		.cost135_12(L135_L[12]),
		.cost135_13(L135_L[13]),
		.cost135_14(L135_L[14]),
		.cost135_15(L135_L[15]),
		.cost135_16(L135_L[16]),
		.cost135_17(L135_L[17]),
		.cost135_18(L135_L[18]),
		.cost135_19(L135_L[19]),
		.cost135_20(L135_L[20]),
		.cost135_21(L135_L[21]),
		.cost135_22(L135_L[22]),
		.cost135_23(L135_L[23]),
		.cost135_24(L135_L[24]),
		.cost135_25(L135_L[25]),
		.cost135_26(L135_L[26]),
		.cost135_27(L135_L[27]),
		.cost135_28(L135_L[28]),
		.cost135_29(L135_L[29]),
		.cost135_30(L135_L[30]),
		.cost135_31(L135_L[31]),
		.cost135_32(L135_L[32]),
		.cost135_33(L135_L[33]),
		.cost135_34(L135_L[34]),
		.cost135_35(L135_L[35]),
		.cost135_36(L135_L[36]),
		.cost135_37(L135_L[37]),
		.cost135_38(L135_L[38]),
		.cost135_39(L135_L[39]),
		.cost135_40(L135_L[40]),
		.cost135_41(L135_L[41]),
		.cost135_42(L135_L[42]),
		.cost135_43(L135_L[43]),
		.cost135_44(L135_L[44]),
		.cost135_45(L135_L[45]),
		.cost135_46(L135_L[46]),
		.cost135_47(L135_L[47]),
		.cost135_48(L135_L[48]),
		.cost135_49(L135_L[49]),
		.cost135_50(L135_L[50]),
		.cost135_51(L135_L[51]),
		.cost135_52(L135_L[52]),
		.cost135_53(L135_L[53]),
		.cost135_54(L135_L[54]),
		.cost135_55(L135_L[55]),
		.cost135_56(L135_L[56]),
		.cost135_57(L135_L[57]),
		.cost135_58(L135_L[58]),
		.cost135_59(L135_L[59]),
		.cost135_60(L135_L[60]),
		.cost135_61(L135_L[61]),
		.cost135_62(L135_L[62]),
		.cost135_63(L135_L[63]),
		
		.L0_0(L_2_0_L[0]),
		.L0_1(L_2_0_L[1]),
		.L0_2(L_2_0_L[2]),
		.L0_3(L_2_0_L[3]),
		.L0_4(L_2_0_L[4]),
		.L0_5(L_2_0_L[5]),
		.L0_6(L_2_0_L[6]),
		.L0_7(L_2_0_L[7]),
		.L0_8(L_2_0_L[8]),
		.L0_9(L_2_0_L[9]),
		.L0_10(L_2_0_L[10]),
		.L0_11(L_2_0_L[11]),
		.L0_12(L_2_0_L[12]),
		.L0_13(L_2_0_L[13]),
		.L0_14(L_2_0_L[14]),
		.L0_15(L_2_0_L[15]),
		.L0_16(L_2_0_L[16]),
		.L0_17(L_2_0_L[17]),
		.L0_18(L_2_0_L[18]),
		.L0_19(L_2_0_L[19]),
		.L0_20(L_2_0_L[20]),
		.L0_21(L_2_0_L[21]),
		.L0_22(L_2_0_L[22]),
		.L0_23(L_2_0_L[23]),
		.L0_24(L_2_0_L[24]),
		.L0_25(L_2_0_L[25]),
		.L0_26(L_2_0_L[26]),
		.L0_27(L_2_0_L[27]),
		.L0_28(L_2_0_L[28]),
		.L0_29(L_2_0_L[29]),
		.L0_30(L_2_0_L[30]),
		.L0_31(L_2_0_L[31]),
		.L0_32(L_2_0_L[32]),
		.L0_33(L_2_0_L[33]),
		.L0_34(L_2_0_L[34]),
		.L0_35(L_2_0_L[35]),
		.L0_36(L_2_0_L[36]),
		.L0_37(L_2_0_L[37]),
		.L0_38(L_2_0_L[38]),
		.L0_39(L_2_0_L[39]),
		.L0_40(L_2_0_L[40]),
		.L0_41(L_2_0_L[41]),
		.L0_42(L_2_0_L[42]),
		.L0_43(L_2_0_L[43]),
		.L0_44(L_2_0_L[44]),
		.L0_45(L_2_0_L[45]),
		.L0_46(L_2_0_L[46]),
		.L0_47(L_2_0_L[47]),
		.L0_48(L_2_0_L[48]),
		.L0_49(L_2_0_L[49]),
		.L0_50(L_2_0_L[50]),
		.L0_51(L_2_0_L[51]),
		.L0_52(L_2_0_L[52]),
		.L0_53(L_2_0_L[53]),
		.L0_54(L_2_0_L[54]),
		.L0_55(L_2_0_L[55]),
		.L0_56(L_2_0_L[56]),
		.L0_57(L_2_0_L[57]),
		.L0_58(L_2_0_L[58]),
		.L0_59(L_2_0_L[59]),
		.L0_60(L_2_0_L[60]),
		.L0_61(L_2_0_L[61]),
		.L0_62(L_2_0_L[62]),
		.L0_63(L_2_0_L[63]),
		
		
		.L135_0(L_2_135_L[0]),
		.L135_1(L_2_135_L[1]),
		.L135_2(L_2_135_L[2]),
		.L135_3(L_2_135_L[3]),
		.L135_4(L_2_135_L[4]),
		.L135_5(L_2_135_L[5]),
		.L135_6(L_2_135_L[6]),
		.L135_7(L_2_135_L[7]),
		.L135_8(L_2_135_L[8]),
		.L135_9(L_2_135_L[9]),
		.L135_10(L_2_135_L[10]),
		.L135_11(L_2_135_L[11]),
		.L135_12(L_2_135_L[12]),
		.L135_13(L_2_135_L[13]),
		.L135_14(L_2_135_L[14]),
		.L135_15(L_2_135_L[15]),
		.L135_16(L_2_135_L[16]),
		.L135_17(L_2_135_L[17]),
		.L135_18(L_2_135_L[18]),
		.L135_19(L_2_135_L[19]),
		.L135_20(L_2_135_L[20]),
		.L135_21(L_2_135_L[21]),
		.L135_22(L_2_135_L[22]),
		.L135_23(L_2_135_L[23]),
		.L135_24(L_2_135_L[24]),
		.L135_25(L_2_135_L[25]),
		.L135_26(L_2_135_L[26]),
		.L135_27(L_2_135_L[27]),
		.L135_28(L_2_135_L[28]),
		.L135_29(L_2_135_L[29]),
		.L135_30(L_2_135_L[30]),
		.L135_31(L_2_135_L[31]),
		.L135_32(L_2_135_L[32]),
		.L135_33(L_2_135_L[33]),
		.L135_34(L_2_135_L[34]),
		.L135_35(L_2_135_L[35]),
		.L135_36(L_2_135_L[36]),
		.L135_37(L_2_135_L[37]),
		.L135_38(L_2_135_L[38]),
		.L135_39(L_2_135_L[39]),
		.L135_40(L_2_135_L[40]),
		.L135_41(L_2_135_L[41]),
		.L135_42(L_2_135_L[42]),
		.L135_43(L_2_135_L[43]),
		.L135_44(L_2_135_L[44]),
		.L135_45(L_2_135_L[45]),
		.L135_46(L_2_135_L[46]),
		.L135_47(L_2_135_L[47]),
		.L135_48(L_2_135_L[48]),
		.L135_49(L_2_135_L[49]),
		.L135_50(L_2_135_L[50]),
		.L135_51(L_2_135_L[51]),
		.L135_52(L_2_135_L[52]),
		.L135_53(L_2_135_L[53]),
		.L135_54(L_2_135_L[54]),
		.L135_55(L_2_135_L[55]),
		.L135_56(L_2_135_L[56]),
		.L135_57(L_2_135_L[57]),
		.L135_58(L_2_135_L[58]),
		.L135_59(L_2_135_L[59]),
		.L135_60(L_2_135_L[60]),
		.L135_61(L_2_135_L[61]),
		.L135_62(L_2_135_L[62]),
		.L135_63(L_2_135_L[63])
		);
	
	
	third_agg#(cost_width) third_agg_Left(
		.clk(clk),
		.rst(rst),
		.clken(clken0),
		.change(change_L),
		.valid_2(valid_2_L),
		.valid_3(valid_3_L),
		.cost0_0(L_2_0_L[0]),
		.cost0_1(L_2_0_L[1]),
		.cost0_2(L_2_0_L[2]),
		.cost0_3(L_2_0_L[3]),
		.cost0_4(L_2_0_L[4]),
		.cost0_5(L_2_0_L[5]),
		.cost0_6(L_2_0_L[6]),
		.cost0_7(L_2_0_L[7]),
		.cost0_8(L_2_0_L[8]),
		.cost0_9(L_2_0_L[9]),
		.cost0_10(L_2_0_L[10]),
		.cost0_11(L_2_0_L[11]),
		.cost0_12(L_2_0_L[12]),
		.cost0_13(L_2_0_L[13]),
		.cost0_14(L_2_0_L[14]),
		.cost0_15(L_2_0_L[15]),
		.cost0_16(L_2_0_L[16]),
		.cost0_17(L_2_0_L[17]),
		.cost0_18(L_2_0_L[18]),
		.cost0_19(L_2_0_L[19]),
		.cost0_20(L_2_0_L[20]),
		.cost0_21(L_2_0_L[21]),
		.cost0_22(L_2_0_L[22]),
		.cost0_23(L_2_0_L[23]),
		.cost0_24(L_2_0_L[24]),
		.cost0_25(L_2_0_L[25]),
		.cost0_26(L_2_0_L[26]),
		.cost0_27(L_2_0_L[27]),
		.cost0_28(L_2_0_L[28]),
		.cost0_29(L_2_0_L[29]),
		.cost0_30(L_2_0_L[30]),
		.cost0_31(L_2_0_L[31]),
		.cost0_32(L_2_0_L[32]),
		.cost0_33(L_2_0_L[33]),
		.cost0_34(L_2_0_L[34]),
		.cost0_35(L_2_0_L[35]),
		.cost0_36(L_2_0_L[36]),
		.cost0_37(L_2_0_L[37]),
		.cost0_38(L_2_0_L[38]),
		.cost0_39(L_2_0_L[39]),
		.cost0_40(L_2_0_L[40]),
		.cost0_41(L_2_0_L[41]),
		.cost0_42(L_2_0_L[42]),
		.cost0_43(L_2_0_L[43]),
		.cost0_44(L_2_0_L[44]),
		.cost0_45(L_2_0_L[45]),
		.cost0_46(L_2_0_L[46]),
		.cost0_47(L_2_0_L[47]),
		.cost0_48(L_2_0_L[48]),
		.cost0_49(L_2_0_L[49]),
		.cost0_50(L_2_0_L[50]),
		.cost0_51(L_2_0_L[51]),
		.cost0_52(L_2_0_L[52]),
		.cost0_53(L_2_0_L[53]),
		.cost0_54(L_2_0_L[54]),
		.cost0_55(L_2_0_L[55]),
		.cost0_56(L_2_0_L[56]),
		.cost0_57(L_2_0_L[57]),
		.cost0_58(L_2_0_L[58]),
		.cost0_59(L_2_0_L[59]),
		.cost0_60(L_2_0_L[60]),
		.cost0_61(L_2_0_L[61]),
		.cost0_62(L_2_0_L[62]),
		.cost0_63(L_2_0_L[63]),
		
		.cost135_0(L_2_135_L[0]),
		.cost135_1(L_2_135_L[1]),
		.cost135_2(L_2_135_L[2]),
		.cost135_3(L_2_135_L[3]),
		.cost135_4(L_2_135_L[4]),
		.cost135_5(L_2_135_L[5]),
		.cost135_6(L_2_135_L[6]),
		.cost135_7(L_2_135_L[7]),
		.cost135_8(L_2_135_L[8]),
		.cost135_9(L_2_135_L[9]),
		.cost135_10(L_2_135_L[10]),
		.cost135_11(L_2_135_L[11]),
		.cost135_12(L_2_135_L[12]),
		.cost135_13(L_2_135_L[13]),
		.cost135_14(L_2_135_L[14]),
		.cost135_15(L_2_135_L[15]),
		.cost135_16(L_2_135_L[16]),
		.cost135_17(L_2_135_L[17]),
		.cost135_18(L_2_135_L[18]),
		.cost135_19(L_2_135_L[19]),
		.cost135_20(L_2_135_L[20]),
		.cost135_21(L_2_135_L[21]),
		.cost135_22(L_2_135_L[22]),
		.cost135_23(L_2_135_L[23]),
		.cost135_24(L_2_135_L[24]),
		.cost135_25(L_2_135_L[25]),
		.cost135_26(L_2_135_L[26]),
		.cost135_27(L_2_135_L[27]),
		.cost135_28(L_2_135_L[28]),
		.cost135_29(L_2_135_L[29]),
		.cost135_30(L_2_135_L[30]),
		.cost135_31(L_2_135_L[31]),
		.cost135_32(L_2_135_L[32]),
		.cost135_33(L_2_135_L[33]),
		.cost135_34(L_2_135_L[34]),
		.cost135_35(L_2_135_L[35]),
		.cost135_36(L_2_135_L[36]),
		.cost135_37(L_2_135_L[37]),
		.cost135_38(L_2_135_L[38]),
		.cost135_39(L_2_135_L[39]),
		.cost135_40(L_2_135_L[40]),
		.cost135_41(L_2_135_L[41]),
		.cost135_42(L_2_135_L[42]),
		.cost135_43(L_2_135_L[43]),
		.cost135_44(L_2_135_L[44]),
		.cost135_45(L_2_135_L[45]),
		.cost135_46(L_2_135_L[46]),
		.cost135_47(L_2_135_L[47]),
		.cost135_48(L_2_135_L[48]),
		.cost135_49(L_2_135_L[49]),
		.cost135_50(L_2_135_L[50]),
		.cost135_51(L_2_135_L[51]),
		.cost135_52(L_2_135_L[52]),
		.cost135_53(L_2_135_L[53]),
		.cost135_54(L_2_135_L[54]),
		.cost135_55(L_2_135_L[55]),
		.cost135_56(L_2_135_L[56]),
		.cost135_57(L_2_135_L[57]),
		.cost135_58(L_2_135_L[58]),
		.cost135_59(L_2_135_L[59]),
		.cost135_60(L_2_135_L[60]),
		.cost135_61(L_2_135_L[61]),
		.cost135_62(L_2_135_L[62]),
		.cost135_63(L_2_135_L[63]),
		
		.agg3_0_0(new3_L0_L[0]),
		.agg3_0_1(new3_L0_L[1]),
		.agg3_0_2(new3_L0_L[2]),
		.agg3_0_3(new3_L0_L[3]),
		.agg3_0_4(new3_L0_L[4]),
		.agg3_0_5(new3_L0_L[5]),
		.agg3_0_6(new3_L0_L[6]),
		.agg3_0_7(new3_L0_L[7]),
		.agg3_0_8(new3_L0_L[8]),
		.agg3_0_9(new3_L0_L[9]),
		.agg3_0_10(new3_L0_L[10]),
		.agg3_0_11(new3_L0_L[11]),
		.agg3_0_12(new3_L0_L[12]),
		.agg3_0_13(new3_L0_L[13]),
		.agg3_0_14(new3_L0_L[14]),
		.agg3_0_15(new3_L0_L[15]),
		.agg3_0_16(new3_L0_L[16]),
		.agg3_0_17(new3_L0_L[17]),
		.agg3_0_18(new3_L0_L[18]),
		.agg3_0_19(new3_L0_L[19]),
		.agg3_0_20(new3_L0_L[20]),
		.agg3_0_21(new3_L0_L[21]),
		.agg3_0_22(new3_L0_L[22]),
		.agg3_0_23(new3_L0_L[23]),
		.agg3_0_24(new3_L0_L[24]),
		.agg3_0_25(new3_L0_L[25]),
		.agg3_0_26(new3_L0_L[26]),
		.agg3_0_27(new3_L0_L[27]),
		.agg3_0_28(new3_L0_L[28]),
		.agg3_0_29(new3_L0_L[29]),
		.agg3_0_30(new3_L0_L[30]),
		.agg3_0_31(new3_L0_L[31]),
		.agg3_0_32(new3_L0_L[32]),
		.agg3_0_33(new3_L0_L[33]),
		.agg3_0_34(new3_L0_L[34]),
		.agg3_0_35(new3_L0_L[35]),
		.agg3_0_36(new3_L0_L[36]),
		.agg3_0_37(new3_L0_L[37]),
		.agg3_0_38(new3_L0_L[38]),
		.agg3_0_39(new3_L0_L[39]),
		.agg3_0_40(new3_L0_L[40]),
		.agg3_0_41(new3_L0_L[41]),
		.agg3_0_42(new3_L0_L[42]),
		.agg3_0_43(new3_L0_L[43]),
		.agg3_0_44(new3_L0_L[44]),
		.agg3_0_45(new3_L0_L[45]),
		.agg3_0_46(new3_L0_L[46]),
		.agg3_0_47(new3_L0_L[47]),
		.agg3_0_48(new3_L0_L[48]),
		.agg3_0_49(new3_L0_L[49]),
		.agg3_0_50(new3_L0_L[50]),
		.agg3_0_51(new3_L0_L[51]),
		.agg3_0_52(new3_L0_L[52]),
		.agg3_0_53(new3_L0_L[53]),
		.agg3_0_54(new3_L0_L[54]),
		.agg3_0_55(new3_L0_L[55]),
		.agg3_0_56(new3_L0_L[56]),
		.agg3_0_57(new3_L0_L[57]),
		.agg3_0_58(new3_L0_L[58]),
		.agg3_0_59(new3_L0_L[59]),
		.agg3_0_60(new3_L0_L[60]),
		.agg3_0_61(new3_L0_L[61]),
		.agg3_0_62(new3_L0_L[62]),
		.agg3_0_63(new3_L0_L[63]),
	
		.agg3_135_0(new3_L135_L[0]),
		.agg3_135_1(new3_L135_L[1]),
		.agg3_135_2(new3_L135_L[2]),
		.agg3_135_3(new3_L135_L[3]),
		.agg3_135_4(new3_L135_L[4]),
		.agg3_135_5(new3_L135_L[5]),
		.agg3_135_6(new3_L135_L[6]),
		.agg3_135_7(new3_L135_L[7]),
		.agg3_135_8(new3_L135_L[8]),
		.agg3_135_9(new3_L135_L[9]),
		.agg3_135_10(new3_L135_L[10]),
		.agg3_135_11(new3_L135_L[11]),
		.agg3_135_12(new3_L135_L[12]),
		.agg3_135_13(new3_L135_L[13]),
		.agg3_135_14(new3_L135_L[14]),
		.agg3_135_15(new3_L135_L[15]),
		.agg3_135_16(new3_L135_L[16]),
		.agg3_135_17(new3_L135_L[17]),
		.agg3_135_18(new3_L135_L[18]),
		.agg3_135_19(new3_L135_L[19]),
		.agg3_135_20(new3_L135_L[20]),
		.agg3_135_21(new3_L135_L[21]),
		.agg3_135_22(new3_L135_L[22]),
		.agg3_135_23(new3_L135_L[23]),
		.agg3_135_24(new3_L135_L[24]),
		.agg3_135_25(new3_L135_L[25]),
		.agg3_135_26(new3_L135_L[26]),
		.agg3_135_27(new3_L135_L[27]),
		.agg3_135_28(new3_L135_L[28]),
		.agg3_135_29(new3_L135_L[29]),
		.agg3_135_30(new3_L135_L[30]),
		.agg3_135_31(new3_L135_L[31]),
		.agg3_135_32(new3_L135_L[32]),
		.agg3_135_33(new3_L135_L[33]),
		.agg3_135_34(new3_L135_L[34]),
		.agg3_135_35(new3_L135_L[35]),
		.agg3_135_36(new3_L135_L[36]),
		.agg3_135_37(new3_L135_L[37]),
		.agg3_135_38(new3_L135_L[38]),
		.agg3_135_39(new3_L135_L[39]),
		.agg3_135_40(new3_L135_L[40]),
		.agg3_135_41(new3_L135_L[41]),
		.agg3_135_42(new3_L135_L[42]),
		.agg3_135_43(new3_L135_L[43]),
		.agg3_135_44(new3_L135_L[44]),
		.agg3_135_45(new3_L135_L[45]),
		.agg3_135_46(new3_L135_L[46]),
		.agg3_135_47(new3_L135_L[47]),
		.agg3_135_48(new3_L135_L[48]),
		.agg3_135_49(new3_L135_L[49]),
		.agg3_135_50(new3_L135_L[50]),
		.agg3_135_51(new3_L135_L[51]),
		.agg3_135_52(new3_L135_L[52]),
		.agg3_135_53(new3_L135_L[53]),
		.agg3_135_54(new3_L135_L[54]),
		.agg3_135_55(new3_L135_L[55]),
		.agg3_135_56(new3_L135_L[56]),
		.agg3_135_57(new3_L135_L[57]),
		.agg3_135_58(new3_L135_L[58]),
		.agg3_135_59(new3_L135_L[59]),
		.agg3_135_60(new3_L135_L[60]),
		.agg3_135_61(new3_L135_L[61]),
		.agg3_135_62(new3_L135_L[62]),
		.agg3_135_63(new3_L135_L[63]),
		
		.L0_0(L_3_0_L[0]),
		.L0_1(L_3_0_L[1]),
		.L0_2(L_3_0_L[2]),
		.L0_3(L_3_0_L[3]),
		.L0_4(L_3_0_L[4]),
		.L0_5(L_3_0_L[5]),
		.L0_6(L_3_0_L[6]),
		.L0_7(L_3_0_L[7]),
		.L0_8(L_3_0_L[8]),
		.L0_9(L_3_0_L[9]),
		.L0_10(L_3_0_L[10]),
		.L0_11(L_3_0_L[11]),
		.L0_12(L_3_0_L[12]),
		.L0_13(L_3_0_L[13]),
		.L0_14(L_3_0_L[14]),
		.L0_15(L_3_0_L[15]),
		.L0_16(L_3_0_L[16]),
		.L0_17(L_3_0_L[17]),
		.L0_18(L_3_0_L[18]),
		.L0_19(L_3_0_L[19]),
		.L0_20(L_3_0_L[20]),
		.L0_21(L_3_0_L[21]),
		.L0_22(L_3_0_L[22]),
		.L0_23(L_3_0_L[23]),
		.L0_24(L_3_0_L[24]),
		.L0_25(L_3_0_L[25]),
		.L0_26(L_3_0_L[26]),
		.L0_27(L_3_0_L[27]),
		.L0_28(L_3_0_L[28]),
		.L0_29(L_3_0_L[29]),
		.L0_30(L_3_0_L[30]),
		.L0_31(L_3_0_L[31]),
		.L0_32(L_3_0_L[32]),
		.L0_33(L_3_0_L[33]),
		.L0_34(L_3_0_L[34]),
		.L0_35(L_3_0_L[35]),
		.L0_36(L_3_0_L[36]),
		.L0_37(L_3_0_L[37]),
		.L0_38(L_3_0_L[38]),
		.L0_39(L_3_0_L[39]),
		.L0_40(L_3_0_L[40]),
		.L0_41(L_3_0_L[41]),
		.L0_42(L_3_0_L[42]),
		.L0_43(L_3_0_L[43]),
		.L0_44(L_3_0_L[44]),
		.L0_45(L_3_0_L[45]),
		.L0_46(L_3_0_L[46]),
		.L0_47(L_3_0_L[47]),
		.L0_48(L_3_0_L[48]),
		.L0_49(L_3_0_L[49]),
		.L0_50(L_3_0_L[50]),
		.L0_51(L_3_0_L[51]),
		.L0_52(L_3_0_L[52]),
		.L0_53(L_3_0_L[53]),
		.L0_54(L_3_0_L[54]),
		.L0_55(L_3_0_L[55]),
		.L0_56(L_3_0_L[56]),
		.L0_57(L_3_0_L[57]),
		.L0_58(L_3_0_L[58]),
		.L0_59(L_3_0_L[59]),
		.L0_60(L_3_0_L[60]),
		.L0_61(L_3_0_L[61]),
		.L0_62(L_3_0_L[62]),
		.L0_63(L_3_0_L[63]),
	
		.L135_0(L_3_135_L[0]),
		.L135_1(L_3_135_L[1]),
		.L135_2(L_3_135_L[2]),
		.L135_3(L_3_135_L[3]),
		.L135_4(L_3_135_L[4]),
		.L135_5(L_3_135_L[5]),
		.L135_6(L_3_135_L[6]),
		.L135_7(L_3_135_L[7]),
		.L135_8(L_3_135_L[8]),
		.L135_9(L_3_135_L[9]),
		.L135_10(L_3_135_L[10]),
		.L135_11(L_3_135_L[11]),
		.L135_12(L_3_135_L[12]),
		.L135_13(L_3_135_L[13]),
		.L135_14(L_3_135_L[14]),
		.L135_15(L_3_135_L[15]),
		.L135_16(L_3_135_L[16]),
		.L135_17(L_3_135_L[17]),
		.L135_18(L_3_135_L[18]),
		.L135_19(L_3_135_L[19]),
		.L135_20(L_3_135_L[20]),
		.L135_21(L_3_135_L[21]),
		.L135_22(L_3_135_L[22]),
		.L135_23(L_3_135_L[23]),
		.L135_24(L_3_135_L[24]),
		.L135_25(L_3_135_L[25]),
		.L135_26(L_3_135_L[26]),
		.L135_27(L_3_135_L[27]),
		.L135_28(L_3_135_L[28]),
		.L135_29(L_3_135_L[29]),
		.L135_30(L_3_135_L[30]),
		.L135_31(L_3_135_L[31]),
		.L135_32(L_3_135_L[32]),
		.L135_33(L_3_135_L[33]),
		.L135_34(L_3_135_L[34]),
		.L135_35(L_3_135_L[35]),
		.L135_36(L_3_135_L[36]),
		.L135_37(L_3_135_L[37]),
		.L135_38(L_3_135_L[38]),
		.L135_39(L_3_135_L[39]),
		.L135_40(L_3_135_L[40]),
		.L135_41(L_3_135_L[41]),
		.L135_42(L_3_135_L[42]),
		.L135_43(L_3_135_L[43]),
		.L135_44(L_3_135_L[44]),
		.L135_45(L_3_135_L[45]),
		.L135_46(L_3_135_L[46]),
		.L135_47(L_3_135_L[47]),
		.L135_48(L_3_135_L[48]),
		.L135_49(L_3_135_L[49]),
		.L135_50(L_3_135_L[50]),
		.L135_51(L_3_135_L[51]),
		.L135_52(L_3_135_L[52]),
		.L135_53(L_3_135_L[53]),
		.L135_54(L_3_135_L[54]),
		.L135_55(L_3_135_L[55]),
		.L135_56(L_3_135_L[56]),
		.L135_57(L_3_135_L[57]),
		.L135_58(L_3_135_L[58]),
		.L135_59(L_3_135_L[59]),
		.L135_60(L_3_135_L[60]),
		.L135_61(L_3_135_L[61]),
		.L135_62(L_3_135_L[62]),
		.L135_63(L_3_135_L[63])
		
		);
	
	
		wire [(cost_width*8-1):0] din_0_L_1 = {L_0_L[7][0],L_0_L[6][0],L_0_L[5][0],L_0_L[4][0],L_0_L[3][0],L_0_L[2][0],L_0_L[1][0],L_0_L[0][0]};
		wire [(cost_width*8-1):0] din_0_L_2 = {L_0_L[15][0],L_0_L[14][0],L_0_L[13][0],L_0_L[12][0],L_0_L[11][0],L_0_L[10][0],L_0_L[9][0],L_0_L[8][0]};
		wire [(cost_width*8-1):0] din_0_L_3 = {L_0_L[23][0],L_0_L[22][0],L_0_L[21][0],L_0_L[20][0],L_0_L[19][0],L_0_L[18][0],L_0_L[17][0],L_0_L[16][0]};
		wire [(cost_width*8-1):0] din_0_L_4 = {L_0_L[31][0],L_0_L[30][0],L_0_L[29][0],L_0_L[28][0],L_0_L[27][0],L_0_L[26][0],L_0_L[25][0],L_0_L[24][0]};
		wire [(cost_width*8-1):0] din_0_L_5 = {L_0_L[39][0],L_0_L[38][0],L_0_L[37][0],L_0_L[36][0],L_0_L[35][0],L_0_L[34][0],L_0_L[33][0],L_0_L[32][0]};
		wire [(cost_width*8-1):0] din_0_L_6 = {L_0_L[47][0],L_0_L[46][0],L_0_L[45][0],L_0_L[44][0],L_0_L[43][0],L_0_L[42][0],L_0_L[41][0],L_0_L[40][0]};
		wire [(cost_width*8-1):0] din_0_L_7 = {L_0_L[55][0],L_0_L[54][0],L_0_L[53][0],L_0_L[52][0],L_0_L[51][0],L_0_L[50][0],L_0_L[49][0],L_0_L[48][0]};
		wire [(cost_width*8-1):0] din_0_L_8 = {L_0_L[63][0],L_0_L[62][0],L_0_L[61][0],L_0_L[60][0],L_0_L[59][0],L_0_L[58][0],L_0_L[57][0],L_0_L[56][0]};
		
		wire [(cost_width*64-1):0] din_0_L = {din_0_L_8,din_0_L_7,din_0_L_6,din_0_L_5,din_0_L_4,din_0_L_3,din_0_L_2,din_0_L_1};
		wire [(cost_width*64-1):0] dout_0_L = Q_Aggregation0_Ram_2[(cost_width*128-1):(cost_width*64)];
	
		genvar k;
		generate for(k=0;k<64;k=k+1) begin: loop3
				assign L_0_L[k][1] = dout_0_L[k*cost_width+(cost_width-1):k*cost_width];
			end
		endgenerate
		
		//135
		wire [((cost_width-2)*8-1):0] din_135_L_1 = {L_135_L[7][0],L_135_L[6][0],L_135_L[5][0],L_135_L[4][0],L_135_L[3][0],L_135_L[2][0],L_135_L[1][0],L_135_L[0][0]};
		wire [((cost_width-2)*8-1):0] din_135_L_2 = {L_135_L[15][0],L_135_L[14][0],L_135_L[13][0],L_135_L[12][0],L_135_L[11][0],L_135_L[10][0],L_135_L[9][0],L_135_L[8][0]};
		wire [((cost_width-2)*8-1):0] din_135_L_3 = {L_135_L[23][0],L_135_L[22][0],L_135_L[21][0],L_135_L[20][0],L_135_L[19][0],L_135_L[18][0],L_135_L[17][0],L_135_L[16][0]};
		wire [((cost_width-2)*8-1):0] din_135_L_4 = {L_135_L[31][0],L_135_L[30][0],L_135_L[29][0],L_135_L[28][0],L_135_L[27][0],L_135_L[26][0],L_135_L[25][0],L_135_L[24][0]};
		wire [((cost_width-2)*8-1):0] din_135_L_5 = {L_135_L[39][0],L_135_L[38][0],L_135_L[37][0],L_135_L[36][0],L_135_L[35][0],L_135_L[34][0],L_135_L[33][0],L_135_L[32][0]};
		wire [((cost_width-2)*8-1):0] din_135_L_6 = {L_135_L[47][0],L_135_L[46][0],L_135_L[45][0],L_135_L[44][0],L_135_L[43][0],L_135_L[42][0],L_135_L[41][0],L_135_L[40][0]};
		wire [((cost_width-2)*8-1):0] din_135_L_7 = {L_135_L[55][0],L_135_L[54][0],L_135_L[53][0],L_135_L[52][0],L_135_L[51][0],L_135_L[50][0],L_135_L[49][0],L_135_L[48][0]};
		wire [((cost_width-2)*8-1):0] din_135_L_8 = {L_135_L[63][0],L_135_L[62][0],L_135_L[61][0],L_135_L[60][0],L_135_L[59][0],L_135_L[58][0],L_135_L[57][0],L_135_L[56][0]};
		wire [((cost_width-2)*64-1):0]din_135_L = {din_135_L_8,din_135_L_7,din_135_L_6,din_135_L_5,din_135_L_4,din_135_L_3,din_135_L_2,din_135_L_1};
		wire [((cost_width-2)*64-1):0] dout_135_L = Q_Aggregation135_Ram_2[((cost_width-2)*128-1):((cost_width-2)*64)];
	
		genvar m;
		generate for(m=0;m<64;m=m+1) begin: loop4
				assign L_135_L[m][1] = dout_135_L[m*(cost_width-2)+(cost_width-3):m*(cost_width-2)];
			end
		endgenerate	
	
	
	//Aggregation modules for the right direction		
	agg2#(cost_width) agg2_Left(
		.clk(clk),
		.rst(rst),
		.clken(clken0),
		.en_first(en_first_L_agg2),

        .P1({P1,2'b00}),
        .P2({P2,2'b00}),
		
		.agg0_0(L_0_L[0][2]),
		.agg0_1(L_0_L[1][2]),
		.agg0_2(L_0_L[2][2]),
		.agg0_3(L_0_L[3][2]),
		.agg0_4(L_0_L[4][2]),
		.agg0_5(L_0_L[5][2]),
		.agg0_6(L_0_L[6][2]),
		.agg0_7(L_0_L[7][2]),
		.agg0_8(L_0_L[8][2]),
		.agg0_9(L_0_L[9][2]),
		.agg0_10(L_0_L[10][2]),
		.agg0_11(L_0_L[11][2]),
		.agg0_12(L_0_L[12][2]),
		.agg0_13(L_0_L[13][2]),
		.agg0_14(L_0_L[14][2]),
		.agg0_15(L_0_L[15][2]),
		.agg0_16(L_0_L[16][2]),
		.agg0_17(L_0_L[17][2]),
		.agg0_18(L_0_L[18][2]),
		.agg0_19(L_0_L[19][2]),
		.agg0_20(L_0_L[20][2]),
		.agg0_21(L_0_L[21][2]),
		.agg0_22(L_0_L[22][2]),
		.agg0_23(L_0_L[23][2]),
		.agg0_24(L_0_L[24][2]),
		.agg0_25(L_0_L[25][2]),
		.agg0_26(L_0_L[26][2]),
		.agg0_27(L_0_L[27][2]),
		.agg0_28(L_0_L[28][2]),
		.agg0_29(L_0_L[29][2]),
		.agg0_30(L_0_L[30][2]),
		.agg0_31(L_0_L[31][2]),
		.agg0_32(L_0_L[32][2]),
		.agg0_33(L_0_L[33][2]),
		.agg0_34(L_0_L[34][2]),
		.agg0_35(L_0_L[35][2]),
		.agg0_36(L_0_L[36][2]),
		.agg0_37(L_0_L[37][2]),
		.agg0_38(L_0_L[38][2]),
		.agg0_39(L_0_L[39][2]),
		.agg0_40(L_0_L[40][2]),
		.agg0_41(L_0_L[41][2]),
		.agg0_42(L_0_L[42][2]),
		.agg0_43(L_0_L[43][2]),
		.agg0_44(L_0_L[44][2]),
		.agg0_45(L_0_L[45][2]),
		.agg0_46(L_0_L[46][2]),
		.agg0_47(L_0_L[47][2]),
		.agg0_48(L_0_L[48][2]),
		.agg0_49(L_0_L[49][2]),
		.agg0_50(L_0_L[50][2]),
		.agg0_51(L_0_L[51][2]),
		.agg0_52(L_0_L[52][2]),
		.agg0_53(L_0_L[53][2]),
		.agg0_54(L_0_L[54][2]),
		.agg0_55(L_0_L[55][2]),
		.agg0_56(L_0_L[56][2]),
		.agg0_57(L_0_L[57][2]),
		.agg0_58(L_0_L[58][2]),
		.agg0_59(L_0_L[59][2]),
		.agg0_60(L_0_L[60][2]),
		.agg0_61(L_0_L[61][2]),
		.agg0_62(L_0_L[62][2]),
		.agg0_63(L_0_L[63][2]),
	
		
		.cost0_0(L_0_L[0][1]),
		.cost0_1(L_0_L[1][1]),
		.cost0_2(L_0_L[2][1]),
		.cost0_3(L_0_L[3][1]),
		.cost0_4(L_0_L[4][1]),
		.cost0_5(L_0_L[5][1]),
		.cost0_6(L_0_L[6][1]),
		.cost0_7(L_0_L[7][1]),
		.cost0_8(L_0_L[8][1]),
		.cost0_9(L_0_L[9][1]),
		.cost0_10(L_0_L[10][1]),
		.cost0_11(L_0_L[11][1]),
		.cost0_12(L_0_L[12][1]),
		.cost0_13(L_0_L[13][1]),
		.cost0_14(L_0_L[14][1]),
		.cost0_15(L_0_L[15][1]),
		.cost0_16(L_0_L[16][1]),
		.cost0_17(L_0_L[17][1]),
		.cost0_18(L_0_L[18][1]),
		.cost0_19(L_0_L[19][1]),
		.cost0_20(L_0_L[20][1]),
		.cost0_21(L_0_L[21][1]),
		.cost0_22(L_0_L[22][1]),
		.cost0_23(L_0_L[23][1]),
		.cost0_24(L_0_L[24][1]),
		.cost0_25(L_0_L[25][1]),
		.cost0_26(L_0_L[26][1]),
		.cost0_27(L_0_L[27][1]),
		.cost0_28(L_0_L[28][1]),
		.cost0_29(L_0_L[29][1]),
		.cost0_30(L_0_L[30][1]),
		.cost0_31(L_0_L[31][1]),
		.cost0_32(L_0_L[32][1]),
		.cost0_33(L_0_L[33][1]),
		.cost0_34(L_0_L[34][1]),
		.cost0_35(L_0_L[35][1]),
		.cost0_36(L_0_L[36][1]),
		.cost0_37(L_0_L[37][1]),
		.cost0_38(L_0_L[38][1]),
		.cost0_39(L_0_L[39][1]),
		.cost0_40(L_0_L[40][1]),
		.cost0_41(L_0_L[41][1]),
		.cost0_42(L_0_L[42][1]),
		.cost0_43(L_0_L[43][1]),
		.cost0_44(L_0_L[44][1]),
		.cost0_45(L_0_L[45][1]),
		.cost0_46(L_0_L[46][1]),
		.cost0_47(L_0_L[47][1]),
		.cost0_48(L_0_L[48][1]),
		.cost0_49(L_0_L[49][1]),
		.cost0_50(L_0_L[50][1]),
		.cost0_51(L_0_L[51][1]),
		.cost0_52(L_0_L[52][1]),
		.cost0_53(L_0_L[53][1]),
		.cost0_54(L_0_L[54][1]),
		.cost0_55(L_0_L[55][1]),
		.cost0_56(L_0_L[56][1]),
		.cost0_57(L_0_L[57][1]),
		.cost0_58(L_0_L[58][1]),
		.cost0_59(L_0_L[59][1]),
		.cost0_60(L_0_L[60][1]),
		.cost0_61(L_0_L[61][1]),
		.cost0_62(L_0_L[62][1]),
		.cost0_63(L_0_L[63][1]),
	
		.cost135_0(L_135_L[0][1]),
		.cost135_1(L_135_L[1][1]),
		.cost135_2(L_135_L[2][1]),
		.cost135_3(L_135_L[3][1]),
		.cost135_4(L_135_L[4][1]),
		.cost135_5(L_135_L[5][1]),
		.cost135_6(L_135_L[6][1]),
		.cost135_7(L_135_L[7][1]),
		.cost135_8(L_135_L[8][1]),
		.cost135_9(L_135_L[9][1]),
		.cost135_10(L_135_L[10][1]),
		.cost135_11(L_135_L[11][1]),
		.cost135_12(L_135_L[12][1]),
		.cost135_13(L_135_L[13][1]),
		.cost135_14(L_135_L[14][1]),
		.cost135_15(L_135_L[15][1]),
		.cost135_16(L_135_L[16][1]),
		.cost135_17(L_135_L[17][1]),
		.cost135_18(L_135_L[18][1]),
		.cost135_19(L_135_L[19][1]),
		.cost135_20(L_135_L[20][1]),
		.cost135_21(L_135_L[21][1]),
		.cost135_22(L_135_L[22][1]),
		.cost135_23(L_135_L[23][1]),
		.cost135_24(L_135_L[24][1]),
		.cost135_25(L_135_L[25][1]),
		.cost135_26(L_135_L[26][1]),
		.cost135_27(L_135_L[27][1]),	
		.cost135_28(L_135_L[28][1]),
		.cost135_29(L_135_L[29][1]),
		.cost135_30(L_135_L[30][1]),
		.cost135_31(L_135_L[31][1]),	
		.cost135_32(L_135_L[32][1]),
		.cost135_33(L_135_L[33][1]),
		.cost135_34(L_135_L[34][1]),
		.cost135_35(L_135_L[35][1]),
		.cost135_36(L_135_L[36][1]),
		.cost135_37(L_135_L[37][1]),
		.cost135_38(L_135_L[38][1]),
		.cost135_39(L_135_L[39][1]),
		.cost135_40(L_135_L[40][1]),
		.cost135_41(L_135_L[41][1]),
		.cost135_42(L_135_L[42][1]),
		.cost135_43(L_135_L[43][1]),
		.cost135_44(L_135_L[44][1]),
		.cost135_45(L_135_L[45][1]),
		.cost135_46(L_135_L[46][1]),
		.cost135_47(L_135_L[47][1]),
		.cost135_48(L_135_L[48][1]),
		.cost135_49(L_135_L[49][1]),
		.cost135_50(L_135_L[50][1]),
		.cost135_51(L_135_L[51][1]),
		.cost135_52(L_135_L[52][1]),
		.cost135_53(L_135_L[53][1]),
		.cost135_54(L_135_L[54][1]),
		.cost135_55(L_135_L[55][1]),
		.cost135_56(L_135_L[56][1]),
		.cost135_57(L_135_L[57][1]),
		.cost135_58(L_135_L[58][1]),
		.cost135_59(L_135_L[59][1]),
		.cost135_60(L_135_L[60][1]),
		.cost135_61(L_135_L[61][1]),
		.cost135_62(L_135_L[62][1]),
		.cost135_63(L_135_L[63][1]),
	
		.min_0_in(min_0_L),
		.min_135(min_135_L),
		.min_0_out(min_0_L),
	
		.L0_0(L_0_L[0][2]),
		.L0_1(L_0_L[1][2]),
		.L0_2(L_0_L[2][2]),
		.L0_3(L_0_L[3][2]),
		.L0_4(L_0_L[4][2]),
		.L0_5(L_0_L[5][2]),
		.L0_6(L_0_L[6][2]),
		.L0_7(L_0_L[7][2]),
		.L0_8(L_0_L[8][2]),
		.L0_9(L_0_L[9][2]),
		.L0_10(L_0_L[10][2]),
		.L0_11(L_0_L[11][2]),
		.L0_12(L_0_L[12][2]),
		.L0_13(L_0_L[13][2]),
		.L0_14(L_0_L[14][2]),
		.L0_15(L_0_L[15][2]),
		.L0_16(L_0_L[16][2]),
		.L0_17(L_0_L[17][2]),
		.L0_18(L_0_L[18][2]),
		.L0_19(L_0_L[19][2]),
		.L0_20(L_0_L[20][2]),
		.L0_21(L_0_L[21][2]),
		.L0_22(L_0_L[22][2]),
		.L0_23(L_0_L[23][2]),
		.L0_24(L_0_L[24][2]),
		.L0_25(L_0_L[25][2]),
		.L0_26(L_0_L[26][2]),
		.L0_27(L_0_L[27][2]),
		.L0_28(L_0_L[28][2]),
		.L0_29(L_0_L[29][2]),
		.L0_30(L_0_L[30][2]),
		.L0_31(L_0_L[31][2]),
		.L0_32(L_0_L[32][2]),
		.L0_33(L_0_L[33][2]),
		.L0_34(L_0_L[34][2]),
		.L0_35(L_0_L[35][2]),
		.L0_36(L_0_L[36][2]),
		.L0_37(L_0_L[37][2]),
		.L0_38(L_0_L[38][2]),
		.L0_39(L_0_L[39][2]),
		.L0_40(L_0_L[40][2]),
		.L0_41(L_0_L[41][2]),
		.L0_42(L_0_L[42][2]),
		.L0_43(L_0_L[43][2]),
		.L0_44(L_0_L[44][2]),
		.L0_45(L_0_L[45][2]),
		.L0_46(L_0_L[46][2]),
		.L0_47(L_0_L[47][2]),
		.L0_48(L_0_L[48][2]),
		.L0_49(L_0_L[49][2]),
		.L0_50(L_0_L[50][2]),
		.L0_51(L_0_L[51][2]),
		.L0_52(L_0_L[52][2]),
		.L0_53(L_0_L[53][2]),
		.L0_54(L_0_L[54][2]),
		.L0_55(L_0_L[55][2]),
		.L0_56(L_0_L[56][2]),
		.L0_57(L_0_L[57][2]),
		.L0_58(L_0_L[58][2]),
		.L0_59(L_0_L[59][2]),
		.L0_60(L_0_L[60][2]),
		.L0_61(L_0_L[61][2]),
		.L0_62(L_0_L[62][2]),
		.L0_63(L_0_L[63][2]),
	
		.L135_0(L_135_L[0][2]),
		.L135_1(L_135_L[1][2]),
		.L135_2(L_135_L[2][2]),
		.L135_3(L_135_L[3][2]),
		.L135_4(L_135_L[4][2]),
		.L135_5(L_135_L[5][2]),
		.L135_6(L_135_L[6][2]),
		.L135_7(L_135_L[7][2]),
		.L135_8(L_135_L[8][2]),
		.L135_9(L_135_L[9][2]),
		.L135_10(L_135_L[10][2]),
		.L135_11(L_135_L[11][2]),
		.L135_12(L_135_L[12][2]),
		.L135_13(L_135_L[13][2]),
		.L135_14(L_135_L[14][2]),
		.L135_15(L_135_L[15][2]),
		.L135_16(L_135_L[16][2]),
		.L135_17(L_135_L[17][2]),
		.L135_18(L_135_L[18][2]),
		.L135_19(L_135_L[19][2]),
		.L135_20(L_135_L[20][2]),
		.L135_21(L_135_L[21][2]),
		.L135_22(L_135_L[22][2]),
		.L135_23(L_135_L[23][2]),
		.L135_24(L_135_L[24][2]),
		.L135_25(L_135_L[25][2]),
		.L135_26(L_135_L[26][2]),
		.L135_27(L_135_L[27][2]),	
		.L135_28(L_135_L[28][2]),
		.L135_29(L_135_L[29][2]),
		.L135_30(L_135_L[30][2]),
		.L135_31(L_135_L[31][2]),
		.L135_32(L_135_L[32][2]),
		.L135_33(L_135_L[33][2]),
		.L135_34(L_135_L[34][2]),
		.L135_35(L_135_L[35][2]),
		.L135_36(L_135_L[36][2]),
		.L135_37(L_135_L[37][2]),
		.L135_38(L_135_L[38][2]),
		.L135_39(L_135_L[39][2]),
		.L135_40(L_135_L[40][2]),
		.L135_41(L_135_L[41][2]),
		.L135_42(L_135_L[42][2]),
		.L135_43(L_135_L[43][2]),
		.L135_44(L_135_L[44][2]),
		.L135_45(L_135_L[45][2]),
		.L135_46(L_135_L[46][2]),
		.L135_47(L_135_L[47][2]),
		.L135_48(L_135_L[48][2]),
		.L135_49(L_135_L[49][2]),
		.L135_50(L_135_L[50][2]),
		.L135_51(L_135_L[51][2]),
		.L135_52(L_135_L[52][2]),
		.L135_53(L_135_L[53][2]),
		.L135_54(L_135_L[54][2]),
		.L135_55(L_135_L[55][2]),
		.L135_56(L_135_L[56][2]),
		.L135_57(L_135_L[57][2]),
		.L135_58(L_135_L[58][2]),
		.L135_59(L_135_L[59][2]),
		.L135_60(L_135_L[60][2]),
		.L135_61(L_135_L[61][2]),
		.L135_62(L_135_L[62][2]),
		.L135_63(L_135_L[63][2]),
	
		.cost_valid(cost_valid)
		);
	
	wire [cost_width-1:0] new4_L0_L[63:0];
	wire [cost_width-3:0] new4_L135_L[63:0];
	
	agg4#(cost_width) agg4_Left(
		.clk(clk),
		.rst0(rst0_L),
		.rst(rst),
		.clken(clken0),
		.en_first(en_first_L),//first pixel of every row
		.en_agg4(en_agg4_L),  //when second row comes
	
		.L0_0(cost_L_in[0]),
		.L0_1(cost_L_in[1]),
		.L0_2(cost_L_in[2]),
		.L0_3(cost_L_in[3]),
		.L0_4(cost_L_in[4]),
		.L0_5(cost_L_in[5]),
		.L0_6(cost_L_in[6]),
		.L0_7(cost_L_in[7]),
		.L0_8(cost_L_in[8]),
		.L0_9(cost_L_in[9]),
		.L0_10(cost_L_in[10]),
		.L0_11(cost_L_in[11]),
		.L0_12(cost_L_in[12]),
		.L0_13(cost_L_in[13]),
		.L0_14(cost_L_in[14]),
		.L0_15(cost_L_in[15]),
		.L0_16(cost_L_in[16]),
		.L0_17(cost_L_in[17]),
		.L0_18(cost_L_in[18]),
		.L0_19(cost_L_in[19]),
		.L0_20(cost_L_in[20]),
		.L0_21(cost_L_in[21]),
		.L0_22(cost_L_in[22]),
		.L0_23(cost_L_in[23]),
		.L0_24(cost_L_in[24]),
		.L0_25(cost_L_in[25]),
		.L0_26(cost_L_in[26]),
		.L0_27(cost_L_in[27]),
		.L0_28(cost_L_in[28]),
		.L0_29(cost_L_in[29]),
		.L0_30(cost_L_in[30]),
		.L0_31(cost_L_in[31]),
		.L0_32(cost_L_in[32]),
		.L0_33(cost_L_in[33]),
		.L0_34(cost_L_in[34]),
		.L0_35(cost_L_in[35]),
		.L0_36(cost_L_in[36]),
		.L0_37(cost_L_in[37]),
		.L0_38(cost_L_in[38]),
		.L0_39(cost_L_in[39]),
		.L0_40(cost_L_in[40]),
		.L0_41(cost_L_in[41]),
		.L0_42(cost_L_in[42]),
		.L0_43(cost_L_in[43]),
		.L0_44(cost_L_in[44]),
		.L0_45(cost_L_in[45]),
		.L0_46(cost_L_in[46]),
		.L0_47(cost_L_in[47]),
		.L0_48(cost_L_in[48]),
		.L0_49(cost_L_in[49]),
		.L0_50(cost_L_in[50]),
		.L0_51(cost_L_in[51]),
		.L0_52(cost_L_in[52]),
		.L0_53(cost_L_in[53]),
		.L0_54(cost_L_in[54]),
		.L0_55(cost_L_in[55]),
		.L0_56(cost_L_in[56]),
		.L0_57(cost_L_in[57]),
		.L0_58(cost_L_in[58]),
		.L0_59(cost_L_in[59]),
		.L0_60(cost_L_in[60]),
		.L0_61(cost_L_in[61]),
		.L0_62(cost_L_in[62]),
		.L0_63(cost_L_in[63]),
		
		.L135_0(cost_L_in[0][cost_width-1:2]),
		.L135_1(cost_L_in[1][cost_width-1:2]),
		.L135_2(cost_L_in[2][cost_width-1:2]),
		.L135_3(cost_L_in[3][cost_width-1:2]),
		.L135_4(cost_L_in[4][cost_width-1:2]),
		.L135_5(cost_L_in[5][cost_width-1:2]),
		.L135_6(cost_L_in[6][cost_width-1:2]),
		.L135_7(cost_L_in[7][cost_width-1:2]),
		.L135_8(cost_L_in[8][cost_width-1:2]),
		.L135_9(cost_L_in[9][cost_width-1:2]),
		.L135_10(cost_L_in[10][cost_width-1:2]),
		.L135_11(cost_L_in[11][cost_width-1:2]),
		.L135_12(cost_L_in[12][cost_width-1:2]),
		.L135_13(cost_L_in[13][cost_width-1:2]),
		.L135_14(cost_L_in[14][cost_width-1:2]),
		.L135_15(cost_L_in[15][cost_width-1:2]),
		.L135_16(cost_L_in[16][cost_width-1:2]),
		.L135_17(cost_L_in[17][cost_width-1:2]),
		.L135_18(cost_L_in[18][cost_width-1:2]),
		.L135_19(cost_L_in[19][cost_width-1:2]),
		.L135_20(cost_L_in[20][cost_width-1:2]),
		.L135_21(cost_L_in[21][cost_width-1:2]),
		.L135_22(cost_L_in[22][cost_width-1:2]),
		.L135_23(cost_L_in[23][cost_width-1:2]),
		.L135_24(cost_L_in[24][cost_width-1:2]),
		.L135_25(cost_L_in[25][cost_width-1:2]),
		.L135_26(cost_L_in[26][cost_width-1:2]),
		.L135_27(cost_L_in[27][cost_width-1:2]),
		.L135_28(cost_L_in[28][cost_width-1:2]),
		.L135_29(cost_L_in[29][cost_width-1:2]),
		.L135_30(cost_L_in[30][cost_width-1:2]),
		.L135_31(cost_L_in[31][cost_width-1:2]),
		.L135_32(cost_L_in[32][cost_width-1:2]),
		.L135_33(cost_L_in[33][cost_width-1:2]),
		.L135_34(cost_L_in[34][cost_width-1:2]),
		.L135_35(cost_L_in[35][cost_width-1:2]),
		.L135_36(cost_L_in[36][cost_width-1:2]),
		.L135_37(cost_L_in[37][cost_width-1:2]),
		.L135_38(cost_L_in[38][cost_width-1:2]),
		.L135_39(cost_L_in[39][cost_width-1:2]),
		.L135_40(cost_L_in[40][cost_width-1:2]),
		.L135_41(cost_L_in[41][cost_width-1:2]),
		.L135_42(cost_L_in[42][cost_width-1:2]),
		.L135_43(cost_L_in[43][cost_width-1:2]),
		.L135_44(cost_L_in[44][cost_width-1:2]),
		.L135_45(cost_L_in[45][cost_width-1:2]),
		.L135_46(cost_L_in[46][cost_width-1:2]),
		.L135_47(cost_L_in[47][cost_width-1:2]),
		.L135_48(cost_L_in[48][cost_width-1:2]),
		.L135_49(cost_L_in[49][cost_width-1:2]),
		.L135_50(cost_L_in[50][cost_width-1:2]),
		.L135_51(cost_L_in[51][cost_width-1:2]),
		.L135_52(cost_L_in[52][cost_width-1:2]),
		.L135_53(cost_L_in[53][cost_width-1:2]),
		.L135_54(cost_L_in[54][cost_width-1:2]),
		.L135_55(cost_L_in[55][cost_width-1:2]),
		.L135_56(cost_L_in[56][cost_width-1:2]),
		.L135_57(cost_L_in[57][cost_width-1:2]),
		.L135_58(cost_L_in[58][cost_width-1:2]),
		.L135_59(cost_L_in[59][cost_width-1:2]),
		.L135_60(cost_L_in[60][cost_width-1:2]),
		.L135_61(cost_L_in[61][cost_width-1:2]),
		.L135_62(cost_L_in[62][cost_width-1:2]),
		.L135_63(cost_L_in[63][cost_width-1:2]),
		
		.new_L0_0(new4_L0_L[0]),
		.new_L0_1(new4_L0_L[1]),
		.new_L0_2(new4_L0_L[2]),
		.new_L0_3(new4_L0_L[3]),
		.new_L0_4(new4_L0_L[4]),
		.new_L0_5(new4_L0_L[5]),
		.new_L0_6(new4_L0_L[6]),
		.new_L0_7(new4_L0_L[7]),
		.new_L0_8(new4_L0_L[8]),
		.new_L0_9(new4_L0_L[9]),
		.new_L0_10(new4_L0_L[10]),
		.new_L0_11(new4_L0_L[11]),
		.new_L0_12(new4_L0_L[12]),
		.new_L0_13(new4_L0_L[13]),
		.new_L0_14(new4_L0_L[14]),
		.new_L0_15(new4_L0_L[15]),
		.new_L0_16(new4_L0_L[16]),
		.new_L0_17(new4_L0_L[17]),
		.new_L0_18(new4_L0_L[18]),
		.new_L0_19(new4_L0_L[19]),
		.new_L0_20(new4_L0_L[20]),
		.new_L0_21(new4_L0_L[21]),
		.new_L0_22(new4_L0_L[22]),
		.new_L0_23(new4_L0_L[23]),
		.new_L0_24(new4_L0_L[24]),
		.new_L0_25(new4_L0_L[25]),
		.new_L0_26(new4_L0_L[26]),
		.new_L0_27(new4_L0_L[27]),
		.new_L0_28(new4_L0_L[28]),
		.new_L0_29(new4_L0_L[29]),
		.new_L0_30(new4_L0_L[30]),
		.new_L0_31(new4_L0_L[31]),
		.new_L0_32(new4_L0_L[32]),
		.new_L0_33(new4_L0_L[33]),
		.new_L0_34(new4_L0_L[34]),
		.new_L0_35(new4_L0_L[35]),
		.new_L0_36(new4_L0_L[36]),
		.new_L0_37(new4_L0_L[37]),
		.new_L0_38(new4_L0_L[38]),
		.new_L0_39(new4_L0_L[39]),
		.new_L0_40(new4_L0_L[40]),
		.new_L0_41(new4_L0_L[41]),
		.new_L0_42(new4_L0_L[42]),
		.new_L0_43(new4_L0_L[43]),
		.new_L0_44(new4_L0_L[44]),
		.new_L0_45(new4_L0_L[45]),
		.new_L0_46(new4_L0_L[46]),
		.new_L0_47(new4_L0_L[47]),
		.new_L0_48(new4_L0_L[48]),
		.new_L0_49(new4_L0_L[49]),
		.new_L0_50(new4_L0_L[50]),
		.new_L0_51(new4_L0_L[51]),
		.new_L0_52(new4_L0_L[52]),
		.new_L0_53(new4_L0_L[53]),
		.new_L0_54(new4_L0_L[54]),
		.new_L0_55(new4_L0_L[55]),
		.new_L0_56(new4_L0_L[56]),
		.new_L0_57(new4_L0_L[57]),
		.new_L0_58(new4_L0_L[58]),
		.new_L0_59(new4_L0_L[59]),
		.new_L0_60(new4_L0_L[60]),
		.new_L0_61(new4_L0_L[61]),
		.new_L0_62(new4_L0_L[62]),
		.new_L0_63(new4_L0_L[63]),
		
		.new_L135_0(new4_L135_L[0]),
		.new_L135_1(new4_L135_L[1]),
		.new_L135_2(new4_L135_L[2]),
		.new_L135_3(new4_L135_L[3]),
		.new_L135_4(new4_L135_L[4]),
		.new_L135_5(new4_L135_L[5]),
		.new_L135_6(new4_L135_L[6]),
		.new_L135_7(new4_L135_L[7]),
		.new_L135_8(new4_L135_L[8]),
		.new_L135_9(new4_L135_L[9]),
		.new_L135_10(new4_L135_L[10]),
		.new_L135_11(new4_L135_L[11]),
		.new_L135_12(new4_L135_L[12]),
		.new_L135_13(new4_L135_L[13]),
		.new_L135_14(new4_L135_L[14]),
		.new_L135_15(new4_L135_L[15]),
		.new_L135_16(new4_L135_L[16]),
		.new_L135_17(new4_L135_L[17]),
		.new_L135_18(new4_L135_L[18]),
		.new_L135_19(new4_L135_L[19]),
		.new_L135_20(new4_L135_L[20]),
		.new_L135_21(new4_L135_L[21]),
		.new_L135_22(new4_L135_L[22]),
		.new_L135_23(new4_L135_L[23]),
		.new_L135_24(new4_L135_L[24]),
		.new_L135_25(new4_L135_L[25]),
		.new_L135_26(new4_L135_L[26]),
		.new_L135_27(new4_L135_L[27]),
		.new_L135_28(new4_L135_L[28]),
		.new_L135_29(new4_L135_L[29]),
		.new_L135_30(new4_L135_L[30]),
		.new_L135_31(new4_L135_L[31]),
		.new_L135_32(new4_L135_L[32]),
		.new_L135_33(new4_L135_L[33]),
		.new_L135_34(new4_L135_L[34]),
		.new_L135_35(new4_L135_L[35]),
		.new_L135_36(new4_L135_L[36]),
		.new_L135_37(new4_L135_L[37]),
		.new_L135_38(new4_L135_L[38]),
		.new_L135_39(new4_L135_L[39]),
		.new_L135_40(new4_L135_L[40]),
		.new_L135_41(new4_L135_L[41]),
		.new_L135_42(new4_L135_L[42]),
		.new_L135_43(new4_L135_L[43]),
		.new_L135_44(new4_L135_L[44]),
		.new_L135_45(new4_L135_L[45]),
		.new_L135_46(new4_L135_L[46]),
		.new_L135_47(new4_L135_L[47]),
		.new_L135_48(new4_L135_L[48]),
		.new_L135_49(new4_L135_L[49]),
		.new_L135_50(new4_L135_L[50]),
		.new_L135_51(new4_L135_L[51]),
		.new_L135_52(new4_L135_L[52]),
		.new_L135_53(new4_L135_L[53]),
		.new_L135_54(new4_L135_L[54]),
		.new_L135_55(new4_L135_L[55]),
		.new_L135_56(new4_L135_L[56]),
		.new_L135_57(new4_L135_L[57]),
		.new_L135_58(new4_L135_L[58]),
		.new_L135_59(new4_L135_L[59]),
		.new_L135_60(new4_L135_L[60]),
		.new_L135_61(new4_L135_L[61]),
		.new_L135_62(new4_L135_L[62]),
		.new_L135_63(new4_L135_L[63]),
		.en_agg3(en_agg3_L)
		);
	
	
	
	agg3#(cost_width) agg3_Left(
		.clk(clk),
		.rst0(rst0_L),
		.rst(rst),
		.clken(clken0),
		.en_first(en_first_L),

        .P1(P1),
        .P2(P2),


		.en_agg3(en_agg3_L),
		.L0_0(new4_L0_L[0]),
		.L0_1(new4_L0_L[1]),
		.L0_2(new4_L0_L[2]),
		.L0_3(new4_L0_L[3]),
		.L0_4(new4_L0_L[4]),
		.L0_5(new4_L0_L[5]),
		.L0_6(new4_L0_L[6]),
		.L0_7(new4_L0_L[7]),
		.L0_8(new4_L0_L[8]),
		.L0_9(new4_L0_L[9]),
		.L0_10(new4_L0_L[10]),
		.L0_11(new4_L0_L[11]),
		.L0_12(new4_L0_L[12]),
		.L0_13(new4_L0_L[13]),
		.L0_14(new4_L0_L[14]),
		.L0_15(new4_L0_L[15]),
		.L0_16(new4_L0_L[16]),
		.L0_17(new4_L0_L[17]),
		.L0_18(new4_L0_L[18]),
		.L0_19(new4_L0_L[19]),
		.L0_20(new4_L0_L[20]),
		.L0_21(new4_L0_L[21]),
		.L0_22(new4_L0_L[22]),
		.L0_23(new4_L0_L[23]),
		.L0_24(new4_L0_L[24]),
		.L0_25(new4_L0_L[25]),
		.L0_26(new4_L0_L[26]),
		.L0_27(new4_L0_L[27]),
		.L0_28(new4_L0_L[28]),
		.L0_29(new4_L0_L[29]),
		.L0_30(new4_L0_L[30]),
		.L0_31(new4_L0_L[31]),
		.L0_32(new4_L0_L[32]),
		.L0_33(new4_L0_L[33]),
		.L0_34(new4_L0_L[34]),
		.L0_35(new4_L0_L[35]),
		.L0_36(new4_L0_L[36]),
		.L0_37(new4_L0_L[37]),
		.L0_38(new4_L0_L[38]),
		.L0_39(new4_L0_L[39]),
		.L0_40(new4_L0_L[40]),
		.L0_41(new4_L0_L[41]),
		.L0_42(new4_L0_L[42]),
		.L0_43(new4_L0_L[43]),
		.L0_44(new4_L0_L[44]),
		.L0_45(new4_L0_L[45]),
		.L0_46(new4_L0_L[46]),
		.L0_47(new4_L0_L[47]),
		.L0_48(new4_L0_L[48]),
		.L0_49(new4_L0_L[49]),
		.L0_50(new4_L0_L[50]),
		.L0_51(new4_L0_L[51]),
		.L0_52(new4_L0_L[52]),
		.L0_53(new4_L0_L[53]),
		.L0_54(new4_L0_L[54]),
		.L0_55(new4_L0_L[55]),
		.L0_56(new4_L0_L[56]),
		.L0_57(new4_L0_L[57]),
		.L0_58(new4_L0_L[58]),
		.L0_59(new4_L0_L[59]),
		.L0_60(new4_L0_L[60]),
		.L0_61(new4_L0_L[61]),
		.L0_62(new4_L0_L[62]),
		.L0_63(new4_L0_L[63]),
		
		.L135_0(new4_L135_L[0]),
		.L135_1(new4_L135_L[1]),
		.L135_2(new4_L135_L[2]),
		.L135_3(new4_L135_L[3]),
		.L135_4(new4_L135_L[4]),
		.L135_5(new4_L135_L[5]),
		.L135_6(new4_L135_L[6]),
		.L135_7(new4_L135_L[7]),
		.L135_8(new4_L135_L[8]),
		.L135_9(new4_L135_L[9]),
		.L135_10(new4_L135_L[10]),
		.L135_11(new4_L135_L[11]),
		.L135_12(new4_L135_L[12]),
		.L135_13(new4_L135_L[13]),
		.L135_14(new4_L135_L[14]),
		.L135_15(new4_L135_L[15]),
		.L135_16(new4_L135_L[16]),
		.L135_17(new4_L135_L[17]),
		.L135_18(new4_L135_L[18]),
		.L135_19(new4_L135_L[19]),
		.L135_20(new4_L135_L[20]),
		.L135_21(new4_L135_L[21]),
		.L135_22(new4_L135_L[22]),
		.L135_23(new4_L135_L[23]),
		.L135_24(new4_L135_L[24]),
		.L135_25(new4_L135_L[25]),
		.L135_26(new4_L135_L[26]),
		.L135_27(new4_L135_L[27]),
		.L135_28(new4_L135_L[28]),
		.L135_29(new4_L135_L[29]),
		.L135_30(new4_L135_L[30]),
		.L135_31(new4_L135_L[31]),
		.L135_32(new4_L135_L[32]),
		.L135_33(new4_L135_L[33]),
		.L135_34(new4_L135_L[34]),
		.L135_35(new4_L135_L[35]),
		.L135_36(new4_L135_L[36]),
		.L135_37(new4_L135_L[37]),
		.L135_38(new4_L135_L[38]),
		.L135_39(new4_L135_L[39]),
		.L135_40(new4_L135_L[40]),
		.L135_41(new4_L135_L[41]),
		.L135_42(new4_L135_L[42]),
		.L135_43(new4_L135_L[43]),
		.L135_44(new4_L135_L[44]),
		.L135_45(new4_L135_L[45]),
		.L135_46(new4_L135_L[46]),
		.L135_47(new4_L135_L[47]),
		.L135_48(new4_L135_L[48]),
		.L135_49(new4_L135_L[49]),
		.L135_50(new4_L135_L[50]),
		.L135_51(new4_L135_L[51]),
		.L135_52(new4_L135_L[52]),
		.L135_53(new4_L135_L[53]),
		.L135_54(new4_L135_L[54]),
		.L135_55(new4_L135_L[55]),
		.L135_56(new4_L135_L[56]),
		.L135_57(new4_L135_L[57]),
		.L135_58(new4_L135_L[58]),
		.L135_59(new4_L135_L[59]),
		.L135_60(new4_L135_L[60]),
		.L135_61(new4_L135_L[61]),
		.L135_62(new4_L135_L[62]),
		.L135_63(new4_L135_L[63]),
		
		.min_135(min_135_L),
		.agg135_0(L_135_L[0][2]),
		.agg135_1(L_135_L[1][2]),
		.agg135_2(L_135_L[2][2]),
		.agg135_3(L_135_L[3][2]),
		.agg135_4(L_135_L[4][2]),
		.agg135_5(L_135_L[5][2]),
		.agg135_6(L_135_L[6][2]),
		.agg135_7(L_135_L[7][2]),
		.agg135_8(L_135_L[8][2]),
		.agg135_9(L_135_L[9][2]),
		.agg135_10(L_135_L[10][2]),
		.agg135_11(L_135_L[11][2]),
		.agg135_12(L_135_L[12][2]),
		.agg135_13(L_135_L[13][2]),
		.agg135_14(L_135_L[14][2]),
		.agg135_15(L_135_L[15][2]),
		.agg135_16(L_135_L[16][2]),
		.agg135_17(L_135_L[17][2]),
		.agg135_18(L_135_L[18][2]),
		.agg135_19(L_135_L[19][2]),
		.agg135_20(L_135_L[20][2]),
		.agg135_21(L_135_L[21][2]),
		.agg135_22(L_135_L[22][2]),
		.agg135_23(L_135_L[23][2]),
		.agg135_24(L_135_L[24][2]),
		.agg135_25(L_135_L[25][2]),
		.agg135_26(L_135_L[26][2]),
		.agg135_27(L_135_L[27][2]),
		.agg135_28(L_135_L[28][2]),
		.agg135_29(L_135_L[29][2]),
		.agg135_30(L_135_L[30][2]),
		.agg135_31(L_135_L[31][2]),
		.agg135_32(L_135_L[32][2]),
		.agg135_33(L_135_L[33][2]),
		.agg135_34(L_135_L[34][2]),
		.agg135_35(L_135_L[35][2]),
		.agg135_36(L_135_L[36][2]),
		.agg135_37(L_135_L[37][2]),
		.agg135_38(L_135_L[38][2]),
		.agg135_39(L_135_L[39][2]),
		.agg135_40(L_135_L[40][2]),
		.agg135_41(L_135_L[41][2]),
		.agg135_42(L_135_L[42][2]),
		.agg135_43(L_135_L[43][2]),
		.agg135_44(L_135_L[44][2]),
		.agg135_45(L_135_L[45][2]),
		.agg135_46(L_135_L[46][2]),
		.agg135_47(L_135_L[47][2]),
		.agg135_48(L_135_L[48][2]),
		.agg135_49(L_135_L[49][2]),
		.agg135_50(L_135_L[50][2]),
		.agg135_51(L_135_L[51][2]),
		.agg135_52(L_135_L[52][2]),
		.agg135_53(L_135_L[53][2]),
		.agg135_54(L_135_L[54][2]),
		.agg135_55(L_135_L[55][2]),
		.agg135_56(L_135_L[56][2]),
		.agg135_57(L_135_L[57][2]),
		.agg135_58(L_135_L[58][2]),
		.agg135_59(L_135_L[59][2]),
		.agg135_60(L_135_L[60][2]),
		.agg135_61(L_135_L[61][2]),
		.agg135_62(L_135_L[62][2]),
		.agg135_63(L_135_L[63][2]),
		
		.new_L0_0(new3_L0_L[0]),
		.new_L0_1(new3_L0_L[1]),
		.new_L0_2(new3_L0_L[2]),
		.new_L0_3(new3_L0_L[3]),
		.new_L0_4(new3_L0_L[4]),
		.new_L0_5(new3_L0_L[5]),
		.new_L0_6(new3_L0_L[6]),
		.new_L0_7(new3_L0_L[7]),
		.new_L0_8(new3_L0_L[8]),
		.new_L0_9(new3_L0_L[9]),
		.new_L0_10(new3_L0_L[10]),
		.new_L0_11(new3_L0_L[11]),
		.new_L0_12(new3_L0_L[12]),
		.new_L0_13(new3_L0_L[13]),
		.new_L0_14(new3_L0_L[14]),
		.new_L0_15(new3_L0_L[15]),
		.new_L0_16(new3_L0_L[16]),
		.new_L0_17(new3_L0_L[17]),
		.new_L0_18(new3_L0_L[18]),
		.new_L0_19(new3_L0_L[19]),
		.new_L0_20(new3_L0_L[20]),
		.new_L0_21(new3_L0_L[21]),
		.new_L0_22(new3_L0_L[22]),
		.new_L0_23(new3_L0_L[23]),
		.new_L0_24(new3_L0_L[24]),
		.new_L0_25(new3_L0_L[25]),
		.new_L0_26(new3_L0_L[26]),
		.new_L0_27(new3_L0_L[27]),
		.new_L0_28(new3_L0_L[28]),
		.new_L0_29(new3_L0_L[29]),
		.new_L0_30(new3_L0_L[30]),
		.new_L0_31(new3_L0_L[31]),
		.new_L0_32(new3_L0_L[32]),
		.new_L0_33(new3_L0_L[33]),
		.new_L0_34(new3_L0_L[34]),
		.new_L0_35(new3_L0_L[35]),
		.new_L0_36(new3_L0_L[36]),
		.new_L0_37(new3_L0_L[37]),
		.new_L0_38(new3_L0_L[38]),
		.new_L0_39(new3_L0_L[39]),
		.new_L0_40(new3_L0_L[40]),
		.new_L0_41(new3_L0_L[41]),
		.new_L0_42(new3_L0_L[42]),
		.new_L0_43(new3_L0_L[43]),
		.new_L0_44(new3_L0_L[44]),
		.new_L0_45(new3_L0_L[45]),
		.new_L0_46(new3_L0_L[46]),
		.new_L0_47(new3_L0_L[47]),
		.new_L0_48(new3_L0_L[48]),
		.new_L0_49(new3_L0_L[49]),
		.new_L0_50(new3_L0_L[50]),
		.new_L0_51(new3_L0_L[51]),
		.new_L0_52(new3_L0_L[52]),
		.new_L0_53(new3_L0_L[53]),
		.new_L0_54(new3_L0_L[54]),
		.new_L0_55(new3_L0_L[55]),
		.new_L0_56(new3_L0_L[56]),
		.new_L0_57(new3_L0_L[57]),
		.new_L0_58(new3_L0_L[58]),
		.new_L0_59(new3_L0_L[59]),
		.new_L0_60(new3_L0_L[60]),
		.new_L0_61(new3_L0_L[61]),
		.new_L0_62(new3_L0_L[62]),
		.new_L0_63(new3_L0_L[63]),
		
		.new_L135_0(new3_L135_L[0]),
		.new_L135_1(new3_L135_L[1]),
		.new_L135_2(new3_L135_L[2]),
		.new_L135_3(new3_L135_L[3]),
		.new_L135_4(new3_L135_L[4]),
		.new_L135_5(new3_L135_L[5]),
		.new_L135_6(new3_L135_L[6]),
		.new_L135_7(new3_L135_L[7]),
		.new_L135_8(new3_L135_L[8]),
		.new_L135_9(new3_L135_L[9]),
		.new_L135_10(new3_L135_L[10]),
		.new_L135_11(new3_L135_L[11]),
		.new_L135_12(new3_L135_L[12]),
		.new_L135_13(new3_L135_L[13]),
		.new_L135_14(new3_L135_L[14]),
		.new_L135_15(new3_L135_L[15]),
		.new_L135_16(new3_L135_L[16]),
		.new_L135_17(new3_L135_L[17]),
		.new_L135_18(new3_L135_L[18]),
		.new_L135_19(new3_L135_L[19]),
		.new_L135_20(new3_L135_L[20]),
		.new_L135_21(new3_L135_L[21]),
		.new_L135_22(new3_L135_L[22]),
		.new_L135_23(new3_L135_L[23]),
		.new_L135_24(new3_L135_L[24]),
		.new_L135_25(new3_L135_L[25]),
		.new_L135_26(new3_L135_L[26]),
		.new_L135_27(new3_L135_L[27]),
		.new_L135_28(new3_L135_L[28]),
		.new_L135_29(new3_L135_L[29]),
		.new_L135_30(new3_L135_L[30]),
		.new_L135_31(new3_L135_L[31]),
		.new_L135_32(new3_L135_L[32]),
		.new_L135_33(new3_L135_L[33]),
		.new_L135_34(new3_L135_L[34]),
		.new_L135_35(new3_L135_L[35]),
		.new_L135_36(new3_L135_L[36]),
		.new_L135_37(new3_L135_L[37]),
		.new_L135_38(new3_L135_L[38]),
		.new_L135_39(new3_L135_L[39]),
		.new_L135_40(new3_L135_L[40]),
		.new_L135_41(new3_L135_L[41]),
		.new_L135_42(new3_L135_L[42]),
		.new_L135_43(new3_L135_L[43]),
		.new_L135_44(new3_L135_L[44]),
		.new_L135_45(new3_L135_L[45]),
		.new_L135_46(new3_L135_L[46]),
		.new_L135_47(new3_L135_L[47]),
		.new_L135_48(new3_L135_L[48]),
		.new_L135_49(new3_L135_L[49]),
		.new_L135_50(new3_L135_L[50]),
		.new_L135_51(new3_L135_L[51]),
		.new_L135_52(new3_L135_L[52]),
		.new_L135_53(new3_L135_L[53]),
		.new_L135_54(new3_L135_L[54]),
		.new_L135_55(new3_L135_L[55]),
		.new_L135_56(new3_L135_L[56]),
		.new_L135_57(new3_L135_L[57]),
		.new_L135_58(new3_L135_L[58]),
		.new_L135_59(new3_L135_L[59]),
		.new_L135_60(new3_L135_L[60]),
		.new_L135_61(new3_L135_L[61]),
		.new_L135_62(new3_L135_L[62]),
		.new_L135_63(new3_L135_L[63]),
		.en_disp(en_disp_L),
		.cost_valid(cost_valid)
		);
	//disparity for the right direction
	
	disparity#(cost_width)  disparity_Left(
	
			.rst(rst),
	
			.clk(clk),
	
			.clken(clken0),
	
			.en_disp(en_agg3_L),
	
			//0?
			.aggregateCost0_0(L_0_L[0][2]),
			.aggregateCost0_1(L_0_L[1][2]),
			.aggregateCost0_2(L_0_L[2][2]), 
			.aggregateCost0_3(L_0_L[3][2]),
			.aggregateCost0_4(L_0_L[4][2]),
			.aggregateCost0_5(L_0_L[5][2]), 
			.aggregateCost0_6(L_0_L[6][2]),
			.aggregateCost0_7(L_0_L[7][2]),
			.aggregateCost0_8(L_0_L[8][2]), 
			.aggregateCost0_9(L_0_L[9][2]),
			.aggregateCost0_10(L_0_L[10][2]),
			.aggregateCost0_11(L_0_L[11][2]), 
			.aggregateCost0_12(L_0_L[12][2]),
			.aggregateCost0_13(L_0_L[13][2]),
			.aggregateCost0_14(L_0_L[14][2]), 
			.aggregateCost0_15(L_0_L[15][2]),
			.aggregateCost0_16(L_0_L[16][2]),
			.aggregateCost0_17(L_0_L[17][2]), 
			.aggregateCost0_18(L_0_L[18][2]),
			.aggregateCost0_19(L_0_L[19][2]),
			.aggregateCost0_20(L_0_L[20][2]), 
			.aggregateCost0_21(L_0_L[21][2]),
			.aggregateCost0_22(L_0_L[22][2]),
			.aggregateCost0_23(L_0_L[23][2]), 
			.aggregateCost0_24(L_0_L[24][2]), 
			.aggregateCost0_25(L_0_L[25][2]),
			.aggregateCost0_26(L_0_L[26][2]),
			.aggregateCost0_27(L_0_L[27][2]), 
			.aggregateCost0_28(L_0_L[28][2]), 
			.aggregateCost0_29(L_0_L[29][2]),
			.aggregateCost0_30(L_0_L[30][2]),
			.aggregateCost0_31(L_0_L[31][2]), 
			.aggregateCost0_32(L_0_L[32][2]), 
			.aggregateCost0_33(L_0_L[33][2]),
			.aggregateCost0_34(L_0_L[34][2]),
			.aggregateCost0_35(L_0_L[35][2]), 
			.aggregateCost0_36(L_0_L[36][2]),
			.aggregateCost0_37(L_0_L[37][2]),
			.aggregateCost0_38(L_0_L[38][2]), 
			.aggregateCost0_39(L_0_L[39][2]),
			.aggregateCost0_40(L_0_L[40][2]),
			.aggregateCost0_41(L_0_L[41][2]), 
			.aggregateCost0_42(L_0_L[42][2]),
			.aggregateCost0_43(L_0_L[43][2]),
			.aggregateCost0_44(L_0_L[44][2]), 
			.aggregateCost0_45(L_0_L[45][2]),
			.aggregateCost0_46(L_0_L[46][2]),
			.aggregateCost0_47(L_0_L[47][2]), 
			.aggregateCost0_48(L_0_L[48][2]),
			.aggregateCost0_49(L_0_L[49][2]),
			.aggregateCost0_50(L_0_L[50][2]), 
			.aggregateCost0_51(L_0_L[51][2]),
			.aggregateCost0_52(L_0_L[52][2]),
			.aggregateCost0_53(L_0_L[53][2]), 
			.aggregateCost0_54(L_0_L[54][2]), 
			.aggregateCost0_55(L_0_L[55][2]),
			.aggregateCost0_56(L_0_L[56][2]),
			.aggregateCost0_57(L_0_L[57][2]), 
			.aggregateCost0_58(L_0_L[58][2]), 
			.aggregateCost0_59(L_0_L[59][2]),
			.aggregateCost0_60(L_0_L[60][2]),
			.aggregateCost0_61(L_0_L[61][2]),
			.aggregateCost0_62(L_0_L[62][2]),
			.aggregateCost0_63(L_0_L[63][2]),	
	
			//135?
			.aggregateCost3_0(L_135_L[0][2]),
			.aggregateCost3_1(L_135_L[1][2]),
			.aggregateCost3_2(L_135_L[2][2]), 
			.aggregateCost3_3(L_135_L[3][2]),
			.aggregateCost3_4(L_135_L[4][2]),
			.aggregateCost3_5(L_135_L[5][2]), 
			.aggregateCost3_6(L_135_L[6][2]),
			.aggregateCost3_7(L_135_L[7][2]),
			.aggregateCost3_8(L_135_L[8][2]), 
			.aggregateCost3_9(L_135_L[9][2]),
			.aggregateCost3_10(L_135_L[10][2]),
			.aggregateCost3_11(L_135_L[11][2]), 
			.aggregateCost3_12(L_135_L[12][2]),
			.aggregateCost3_13(L_135_L[13][2]),
			.aggregateCost3_14(L_135_L[14][2]), 
			.aggregateCost3_15(L_135_L[15][2]),
			.aggregateCost3_16(L_135_L[16][2]),
			.aggregateCost3_17(L_135_L[17][2]), 
			.aggregateCost3_18(L_135_L[18][2]),
			.aggregateCost3_19(L_135_L[19][2]),
			.aggregateCost3_20(L_135_L[20][2]), 
			.aggregateCost3_21(L_135_L[21][2]),
			.aggregateCost3_22(L_135_L[22][2]),
			.aggregateCost3_23(L_135_L[23][2]), 
			.aggregateCost3_24(L_135_L[24][2]), 
			.aggregateCost3_25(L_135_L[25][2]),
			.aggregateCost3_26(L_135_L[26][2]),
			.aggregateCost3_27(L_135_L[27][2]), 
			.aggregateCost3_28(L_135_L[28][2]), 
			.aggregateCost3_29(L_135_L[29][2]),
			.aggregateCost3_30(L_135_L[30][2]),
			.aggregateCost3_31(L_135_L[31][2]), 
			.aggregateCost3_32(L_135_L[32][2]), 
			.aggregateCost3_33(L_135_L[33][2]),
			.aggregateCost3_34(L_135_L[34][2]),
			.aggregateCost3_35(L_135_L[35][2]), 
			.aggregateCost3_36(L_135_L[36][2]),
			.aggregateCost3_37(L_135_L[37][2]),
			.aggregateCost3_38(L_135_L[38][2]), 
			.aggregateCost3_39(L_135_L[39][2]),
			.aggregateCost3_40(L_135_L[40][2]),
			.aggregateCost3_41(L_135_L[41][2]), 
			.aggregateCost3_42(L_135_L[42][2]),
			.aggregateCost3_43(L_135_L[43][2]),
			.aggregateCost3_44(L_135_L[44][2]), 
			.aggregateCost3_45(L_135_L[45][2]),
			.aggregateCost3_46(L_135_L[46][2]),
			.aggregateCost3_47(L_135_L[47][2]), 
			.aggregateCost3_48(L_135_L[48][2]),
			.aggregateCost3_49(L_135_L[49][2]),
			.aggregateCost3_50(L_135_L[50][2]), 
			.aggregateCost3_51(L_135_L[51][2]),
			.aggregateCost3_52(L_135_L[52][2]),
			.aggregateCost3_53(L_135_L[53][2]), 
			.aggregateCost3_54(L_135_L[54][2]), 
			.aggregateCost3_55(L_135_L[55][2]),
			.aggregateCost3_56(L_135_L[56][2]),
			.aggregateCost3_57(L_135_L[57][2]), 
			.aggregateCost3_58(L_135_L[58][2]), 
			.aggregateCost3_59(L_135_L[59][2]),
			.aggregateCost3_60(L_135_L[60][2]),
			.aggregateCost3_61(L_135_L[61][2]),
			.aggregateCost3_62(L_135_L[62][2]),
			.aggregateCost3_63(L_135_L[63][2]),
	
			.disp_final(disp_L),
	
			.valid_final(valid_final_L),
	
			.cost_valid(cost_valid)
	
			);
	
	
	
	wire valid_Aggregation0;
	assign D_Aggregation0_Ram_1 = {din_0_L,din_0_R};
	SRAM_control_Aggregation0#((cost_width*128),11,0) SRAM_control_Aggregation0_inst1(
		.clk(clk),
		 .rst(rst),
		.clken(clken0&valid_3_R),
		.width(width-11'd4),
		.wr_en(wr_en_Agg0_inst1),
		.wr_addr(wr_addr_Agg0_inst1),
		.rd_addr(rd_addr_Agg0_inst1),
		.cost_valid(cost_valid),
		.BWEB_s(),
		 .valid()
	);
	//BWEB
    wire[(cost_width*128-1):0] BWEB0;
	assign BWEB0={cost0_valid_B,cost0_valid_B};
//	assign BWEB_Agg0_inst1=wr_en_Agg0_inst1?BWEB0:{(cost_width*128){1'b0}};
	assign BWEB_Agg0_inst1={(cost_width*128){1'b0}};
	wire valid_Aggregation135;
	assign D_Aggregation135_Ram_1 = {din_135_L,din_135_R};

	SRAM_control_Aggregation135#(((cost_width-2)*128),11,0) SRAM_control_Aggregation135_inst1(
		.clk(clk),
		 .rst(rst),
		.clken(clken0&valid_3_R),
		.width(width-11'd4),
		.wr_en(wr_en_Agg135_inst1),
		.wr_addr(wr_addr_Agg135_inst1),
		.rd_addr(rd_addr_Agg135_inst1),
		.cost_valid(cost_valid),
		.BWEB_s(),
		 .valid()
	);
    wire[((cost_width-2)*128-1):0] BWEB135;
	assign BWEB135={cost135_valid_B,cost135_valid_B};
//	assign BWEB_Agg135_inst1=wr_en_Agg135_inst1?BWEB135:{((cost_width-2)*128){1'b0}};
	assign BWEB_Agg135_inst1={((cost_width-2)*128){1'b0}};

	reg [31:0] count;    
	reg [31:0] cnt_first;
	reg [31:0] test;
	wire [31:0] HW ;
	assign HW = width*height;
	always@(posedge clk or negedge rst)begin
		if(rst==0)begin
			count <= 32'd0;
			cnt_first <= 32'd0;
			test <= 32'd0;
			en_agg4_L<=1'd0;
			en_first_L<=1'd0;
			en_first_L_agg2<=1'd0;
			en_agg4_R<=1'd0;
			en_first_R<=1'd0;
			en_first_R_agg2<=1'd0;
			change_L<=1'd0;
			change_R<=1'd0;
			rst0_L<=1'd0;
			rst0_R<=1'd0;
		end
		else if(clken0) begin
			//count<=count+1;
			test<=test+1;
			if(en_L&&en_R)begin
				if(count==HW)begin
					count<=1'd1;
				end
				else begin
					count<=count+1;
				end
				//When the first pixel just come to the input port of Agg4
				if(cnt_first==width-1&&count>=1)begin
					en_first_L<=1'd1;
					en_first_R<=1'd1;
					cnt_first<=1'd1;
				end
				else begin
					en_first_L<=1'd0;
					en_first_R<=1'd0;
					cnt_first<=cnt_first+1;		
				end
				//When the first pixel just come to the input port of Agg2
				if(cnt_first==width-2&&count>=1)begin
					en_first_L_agg2<=1'd1;
					en_first_R_agg2<=1'd1;
				end
				else begin
					en_first_L_agg2<=1'd0;
					en_first_R_agg2<=1'd0;		
				end
				//Change the input data of third agg from second agg to agg3
				if(count>=width+1)begin
					change_L<=1'd1;
					change_R<=1'd1;
				end
				else begin
					change_L<=1'd0;
					change_R<=1'd0;	
				end
				//When the first pixel just come to the input port of Agg4
				if(count>=width-1)begin
					rst0_L<=1'd1;
					rst0_R<=1'd1;
					en_agg4_L<=1'd1;
					en_agg4_R<=1'd1;
				end
				else begin
					rst0_L<=1'd0;
					rst0_R<=1'd0;	
					en_agg4_L<=1'd0;
					en_agg4_R<=1'd0;
				end
			end
		end
	end
	
	endmodule
	
