module LUT_SRT4
(
	//input
	D,
	W,
	//output 
	q1
	
);
	input		[3:0]		D;
	input    [21:0]   W;
	output	[2:0]	q1;
	
	wire [21:0] W_temp1;
	wire [23:0] W_temp2;
        wire [21:0] W_temp3;
	assign W_temp1=W[21]?{1'b1,~W[20:0]+21'd1}:{W};
	//assign W_temp2={W[21],W_temp1[18:0],2'd0};//第一位为符号位//000.00
	assign W_temp2={W_temp1,2'b00};
	assign W_temp3=W[21]?{1'b1,W_temp2[20:0]}:{1'b0,W_temp2[20:0]};
	assign q1=q_temp(W_temp3,D);
	function [2:0] q_temp(input [21:0] W_temp,input [3:0] D);
	case(D)
	4'b1000:q_temp=((W_temp[21]==0) && (W_temp[20:0] >= 21'b00_0011_0000_0000_0000_000))?{3'b010} :
			((W_temp[21]==0) && (21'b00_0001_0000_0000_0000_000 <= W_temp[20:0]) &&( W_temp[20:0] < 21'b00_0011_0000_0000_0000_000))?{3'b001} :
			((W_temp[21]==1) && (W_temp[20:0]>21'b00_0011_0100_0000_0000_000))?{3'b110} :
			((W_temp[21]==1) && (21'b00_0001_0000_0000_0000_000<W_temp[20:0]) && (W_temp[20:0]<=21'b00_0011_0100_0000_0000_000))?{3'b111}:{3'b000};
	4'b1001:q_temp=((W_temp[21]==0) && (W_temp[20:0] >= 21'b00_0011_1000_0000_0000_000))?{3'b010} :
			((W_temp[21]==0) && (21'b00_0001_0000_0000_0000_000 <= W_temp[20:0]) && (W_temp[20:0] < 21'b00_0011_1000_0000_0000_000))?{3'b001} :
			((W_temp[21]==1) && (W_temp[20:0]>21'b00_0011_1000_0000_0000_000))?{3'b110} :
			((W_temp[21]==1) && (21'b00_0001_0000_0000_0000_000 < W_temp[20:0]) && (W_temp[20:0]<=21'b00_0011_1000_0000_0000_000))?{3'b111}:{3'b000};
	4'b1010:q_temp=((W_temp[21]==0) && (W_temp[20:0] >= 21'b00_0011_1100_0000_0000_000))?{3'b010} :
			((W_temp[21]==0) && (21'b00_0001_0000_0000_0000_000 <= W_temp[20:0]) && (W_temp[20:0] < 21'b00_0011_1100_0000_0000_000))?{3'b001} :
			((W_temp[21]==1) && (W_temp[20:0]>21'b00_0100_0000_0000_0000_000))?{3'b110} :
			((W_temp[21]==1) && (21'b00_0001_1000_0000_0000_000 < W_temp[20:0]) && (W_temp[20:0]<=21'b00_0100_0000_0000_0000_000))?{3'b111}:{3'b000};
	4'b1011:q_temp=((W_temp[21]==0) && (W_temp[20:0] >= 21'b00_0100_0000_0000_0000_000))?{3'b010} :
			((W_temp[21]==0) && (21'b00_0001_0000_0000_0000_000 <= W_temp[20:0]) && (W_temp[20:0] < 21'b00_0100_0000_0000_0000_000))?{3'b001} :
			((W_temp[21]==1) && (W_temp[20:0] > 21'b00_0100_1000_0000_0000_000))?{3'b110} :
			((W_temp[21]==1) && (21'b00_0001_1000_0000_0000_000 < W_temp[20:0]<=21'b00_0100_1000_0000_0000_000))?{3'b111}:{3'b000};
	4'b1100:q_temp=((W_temp[21]==0) && (W_temp[20:0] >= 21'b00_0101_0000_0000_0000_000))?{3'b010} :
			((W_temp[21]==0) && (21'b00_0001_1000_0000_0000_000 <= W_temp[20:0]) && (W_temp[20:0] < 21'b00_0101_0000_0000_0000_000))?{3'b001} :
			((W_temp[21]==1) && (W_temp[20:0]>21'b00_0100_1000_0000_0000_000))?{3'b110} :
			((W_temp[21]==1) && (21'b00_0001_1000_0000_0000_000<W_temp[20:0]) && (W_temp[20:0]<=21'b00_0100_1000_0000_0000_000))?{3'b111}:{3'b000};
	4'b1101:q_temp=((W_temp[21]==0) && (W_temp[20:0] >= 21'b00_0100_1100_0000_0000_000))?{3'b010} :
			((W_temp[21]==0) && (21'b00_0001_1000_0000_0000_000 <= W_temp[20:0]) && (W_temp[20:0]  < 21'b00_0100_1100_0000_0000_000))?{3'b001} :
			((W_temp[21]==1) && (W_temp[20:0]>21'b00_0101_0000_0000_0000_000))?{3'b110} :
			((W_temp[21]==1) && (21'b00_0010_0000_0000_0000_000<W_temp[20:0]) && (W_temp[20:0]<=21'b00_0101_0000_0000_0000_000))?{3'b111}:{3'b000};
	4'b1110:q_temp=((W_temp[21]==0) && (W_temp[20:0] >= 21'b00_0101_0000_0000_0000_000))?{3'b010} :
			((W_temp[21]==0) && (21'b00_0010_0000_0000_0000_000 <= W_temp[20:0]) &&(W_temp[20:0] < 21'b00_0101_0000_0000_0000_000))?{3'b001} :
			((W_temp[21]==1) && (W_temp[20:0]>21'b00_0101_1000_0000_0000_000))?{3'b110} :
			((W_temp[21]==1) && (21'b00_0010_0000_0000_0000_000<W_temp[20:0]<=21'b00_0101_1000_0000_0000_000))?{3'b111}:{3'b000};
	4'b1111:q_temp=((W_temp[21]==0) && (W_temp[20:0] >= 21'b00_0110_0000_0000_0000_000))?{3'b010} :
			((W_temp[21]==0) && (21'b00_0010_0000_0000_0000_000 <= W_temp[20:0]) && (W_temp[20:0] < 21'b00_0110_0000_0000_0000_000))?{3'b001} :
			((W_temp[21]==1) && (W_temp[20:0]>21'b00_0110_0000_0000_0000_000))?{3'b110} :
			((W_temp[21]==1) && (21'b00_0010_0000_0000_0000_000 < W_temp[20:0]) && (W_temp[20:0]<=21'b00_0110_0000_0000_0000_000))?{3'b111}:{3'b000};
	default:q_temp=3'b100;
	endcase
endfunction
endmodule
